[
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 3,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            1,
            695
        ],
        "focused": false,
        "bounds": [
            [
                0,
                0
            ],
            [
                1080,
                2400
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.widget.FrameLayout",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": -1,
        "temp_id": 0,
        "size": "1080*2400",
        "signature": "[class]android.widget.FrameLayout[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "bd0083930bf52f52f9c2ee8d3fce09d5",
        "bound_box": "0,0,1080,2400",
        "content_free_signature": "[class]android.widget.FrameLayout[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            2
        ],
        "focused": false,
        "bounds": [
            [
                0,
                0
            ],
            [
                1080,
                2274
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.widget.LinearLayout",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 0,
        "temp_id": 1,
        "size": "1080*2274",
        "signature": "[class]android.widget.LinearLayout[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "6892907490647f5d6911fad9738282e0",
        "bound_box": "0,0,1080,2274",
        "content_free_signature": "[class]android.widget.LinearLayout[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            3
        ],
        "focused": false,
        "bounds": [
            [
                0,
                63
            ],
            [
                1080,
                2274
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.widget.FrameLayout",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 1,
        "temp_id": 2,
        "size": "1080*2211",
        "signature": "[class]android.widget.FrameLayout[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "eb6d4b8ee026b3fa6faf9d020c5cad76",
        "bound_box": "0,63,1080,2274",
        "content_free_signature": "[class]android.widget.FrameLayout[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            4
        ],
        "focused": false,
        "bounds": [
            [
                0,
                63
            ],
            [
                1080,
                2274
            ]
        ],
        "resource_id": "com.android.chrome:id/action_bar_root",
        "checked": false,
        "text": null,
        "class": "android.widget.FrameLayout",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 2,
        "temp_id": 3,
        "size": "1080*2211",
        "signature": "[class]android.widget.FrameLayout[resource_id]com.android.chrome:id/action_bar_root[visible]True[text]None[enabled,,]",
        "view_str": "ee44a51611fbbaca235c29d7be02454b",
        "bound_box": "0,63,1080,2274",
        "content_free_signature": "[class]android.widget.FrameLayout[resource_id]com.android.chrome:id/action_bar_root[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 3,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            5,
            693
        ],
        "focused": false,
        "bounds": [
            [
                0,
                63
            ],
            [
                1080,
                2274
            ]
        ],
        "resource_id": "android:id/content",
        "checked": false,
        "text": null,
        "class": "android.widget.FrameLayout",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 3,
        "temp_id": 4,
        "size": "1080*2211",
        "signature": "[class]android.widget.FrameLayout[resource_id]android:id/content[visible]True[text]None[enabled,,]",
        "view_str": "8f661d0fb75b6b621a5eea75d73d7d34",
        "bound_box": "0,63,1080,2274",
        "content_free_signature": "[class]android.widget.FrameLayout[resource_id]android:id/content[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 3,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            6,
            674
        ],
        "focused": false,
        "bounds": [
            [
                0,
                63
            ],
            [
                1080,
                2274
            ]
        ],
        "resource_id": "com.android.chrome:id/coordinator",
        "checked": false,
        "text": null,
        "class": "android.view.ViewGroup",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 4,
        "temp_id": 5,
        "size": "1080*2211",
        "signature": "[class]android.view.ViewGroup[resource_id]com.android.chrome:id/coordinator[visible]True[text]None[enabled,,]",
        "view_str": "b0b7c8b198f878dbfda08082c1527e3f",
        "bound_box": "0,63,1080,2274",
        "content_free_signature": "[class]android.view.ViewGroup[resource_id]com.android.chrome:id/coordinator[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            7,
            9
        ],
        "focused": false,
        "bounds": [
            [
                0,
                63
            ],
            [
                1080,
                2274
            ]
        ],
        "resource_id": "com.android.chrome:id/compositor_view_holder",
        "checked": false,
        "text": null,
        "class": "android.widget.FrameLayout",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 5,
        "temp_id": 6,
        "size": "1080*2211",
        "signature": "[class]android.widget.FrameLayout[resource_id]com.android.chrome:id/compositor_view_holder[visible]True[text]None[enabled,,]",
        "view_str": "7b765fdfd4bfc523d2bdb44d7f4c01e5",
        "bound_box": "0,63,1080,2274",
        "content_free_signature": "[class]android.widget.FrameLayout[resource_id]com.android.chrome:id/compositor_view_holder[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            8
        ],
        "focused": false,
        "bounds": [
            [
                0,
                63
            ],
            [
                1080,
                2274
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.widget.FrameLayout",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 6,
        "temp_id": 7,
        "size": "1080*2211",
        "signature": "[class]android.widget.FrameLayout[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "1f2a04e5f3ceaa76877afc3376546656",
        "bound_box": "0,63,1080,2274",
        "content_free_signature": "[class]android.widget.FrameLayout[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                63
            ],
            [
                1080,
                2274
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 7,
        "temp_id": 8,
        "size": "1080*2211",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "0039e922c3c52932c64931284a9d0b04",
        "bound_box": "0,63,1080,2274",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            10
        ],
        "focused": false,
        "bounds": [
            [
                0,
                63
            ],
            [
                1080,
                2274
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.widget.FrameLayout",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 6,
        "temp_id": 9,
        "size": "1080*2211",
        "signature": "[class]android.widget.FrameLayout[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "2a020248da6c40f98205da7c21e2fb9e",
        "bound_box": "0,63,1080,2274",
        "content_free_signature": "[class]android.widget.FrameLayout[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [
            11
        ],
        "focused": true,
        "bounds": [
            [
                0,
                210
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "google - Google Search",
        "class": "android.webkit.WebView",
        "scrollable": true,
        "selected": false,
        "long_clickable": false,
        "parent": 9,
        "temp_id": 10,
        "size": "1084*2066",
        "signature": "[class]android.webkit.WebView[resource_id]None[visible]True[text]google - Google Search[enabled,,]",
        "view_str": "31289e2e06a4791c142662ebfd6faa6f",
        "bound_box": "0,210,1084,2276",
        "content_free_signature": "[class]android.webkit.WebView[resource_id]None[visible]True",
        "allowed_actions": [
            "scroll up",
            "scroll down",
            "scroll left",
            "scroll right"
        ],
        "status": [],
        "local_id": "0",
        "full_desc": "<scrollbar bound_box=0,210,1084,2276>google - Google Search</scrollbar>",
        "desc": "<scrollbar bound_box=0,210,1084,2276>google - Google Search</scrollbar>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 8,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            12,
            30,
            31,
            662,
            665
        ],
        "focused": false,
        "bounds": [
            [
                0,
                210
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 10,
        "temp_id": 11,
        "size": "1084*2066",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "94a45214b018e0cb5022ae5d6a98b55c",
        "bound_box": "0,210,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "1",
        "full_desc": "<button bound_box=0,210,1084,2276></button>",
        "desc": "<button bound_box=0,210,1084,2276></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            13,
            19
        ],
        "focused": false,
        "bounds": [
            [
                0,
                210
            ],
            [
                1084,
                519
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 11,
        "temp_id": 12,
        "size": "1084*309",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "82e69468164c9429f58477e81105f192",
        "bound_box": "0,210,1084,519",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            14,
            16
        ],
        "focused": false,
        "bounds": [
            [
                0,
                210
            ],
            [
                1084,
                378
            ]
        ],
        "resource_id": "qslc",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 12,
        "temp_id": 13,
        "size": "1084*168",
        "signature": "[class]android.view.View[resource_id]qslc[visible]True[text][enabled,,]",
        "view_str": "85309c44f4029d0be22e29641d47c817",
        "bound_box": "0,210,1084,378",
        "content_free_signature": "[class]android.view.View[resource_id]qslc[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google",
        "children": [
            15
        ],
        "focused": false,
        "bounds": [
            [
                420,
                210
            ],
            [
                664,
                393
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 13,
        "temp_id": 14,
        "size": "244*183",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "dd9a610eff4a510d9ebbfe506d2e2e08",
        "bound_box": "420,210,664,393",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "2",
        "full_desc": "<button alt='Google' bound_box=420,210,664,393></button>",
        "desc": "<button alt='Google' bound_box=420,210,664,393></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                420,
                252
            ],
            [
                664,
                349
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "This image isn‘t labeled. Open the More Options menu at the top right to get image descriptions.",
        "class": "android.widget.Image",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 14,
        "temp_id": 15,
        "size": "244*97",
        "signature": "[class]android.widget.Image[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "28620763e400da96b9b81ca5cbcb92ff",
        "bound_box": "420,252,664,349",
        "content_free_signature": "[class]android.widget.Image[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "3",
        "full_desc": "<button bound_box=420,252,664,349>This image isn‘t labeled. Open the More Options me</button>",
        "desc": "<button bound_box=420,252,664,349>This image isn‘t labeled. Open the More Options me</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            17
        ],
        "focused": false,
        "bounds": [
            [
                913,
                210
            ],
            [
                1084,
                370
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 13,
        "temp_id": 16,
        "size": "171*160",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "cededc43922d5a989cd0508e7f3dc1a3",
        "bound_box": "913,210,1084,370",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [
            18
        ],
        "focused": false,
        "bounds": [
            [
                945,
                217
            ],
            [
                1073,
                349
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google Account: Agent Test (testmobileagent11@gmail.com)",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 16,
        "temp_id": 17,
        "size": "128*132",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "1c079a270a25349a0549d3e9d5588223",
        "bound_box": "945,217,1073,349",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "4",
        "full_desc": "<button bound_box=945,217,1073,349>Google Account: Agent Test (testmobileagent11@gmai</button>",
        "desc": "<button bound_box=945,217,1073,349>Google Account: Agent Test (testmobileagent11@gmai</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                955,
                231
            ],
            [
                1063,
                336
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google Account: Agent Test (testmobileagent11@gmail.com)",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 17,
        "temp_id": 18,
        "size": "108*105",
        "signature": "[class]android.widget.Button[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "a5ca28ed117b09ef67fe18d4906eaf75",
        "bound_box": "955,231,1063,336",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "5",
        "full_desc": "<button bound_box=955,231,1063,336>Google Account: Agent Test (testmobileagent11@gmai</button>",
        "desc": "<button bound_box=955,231,1063,336>Google Account: Agent Test (testmobileagent11@gmai</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            20
        ],
        "focused": false,
        "bounds": [
            [
                42,
                372
            ],
            [
                1042,
                493
            ]
        ],
        "resource_id": "sfcnt",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 12,
        "temp_id": 19,
        "size": "1000*121",
        "signature": "[class]android.view.View[resource_id]sfcnt[visible]True[text][enabled,,]",
        "view_str": "811ce77671af073b3dff6ed645778f6f",
        "bound_box": "42,372,1042,493",
        "content_free_signature": "[class]android.view.View[resource_id]sfcnt[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            21
        ],
        "focused": false,
        "bounds": [
            [
                42,
                372
            ],
            [
                1042,
                493
            ]
        ],
        "resource_id": "gws-quantum-experimental_page_header__sbox",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 19,
        "temp_id": 20,
        "size": "1000*121",
        "signature": "[class]android.view.View[resource_id]gws-quantum-experimental_page_header__sbox[visible]True[text][enabled,,]",
        "view_str": "166c588df108e8af74569faf619f86c0",
        "bound_box": "42,372,1042,493",
        "content_free_signature": "[class]android.view.View[resource_id]gws-quantum-experimental_page_header__sbox[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 7,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            22,
            23,
            24,
            26,
            27,
            28
        ],
        "focused": false,
        "bounds": [
            [
                42,
                372
            ],
            [
                1042,
                493
            ]
        ],
        "resource_id": "tsf",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 20,
        "temp_id": 21,
        "size": "1000*121",
        "signature": "[class]android.view.View[resource_id]tsf[visible]True[text][enabled,,]",
        "view_str": "0d4de5017125c7112127cb4312b5a207",
        "bound_box": "42,372,1042,493",
        "content_free_signature": "[class]android.view.View[resource_id]tsf[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                372
            ],
            [
                1042,
                504
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 21,
        "temp_id": 22,
        "size": "1000*132",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "319dc4c1fce8d2135fa87d7a336ce880",
        "bound_box": "42,372,1042,504",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                372
            ],
            [
                168,
                493
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google Search",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 21,
        "temp_id": 23,
        "size": "126*121",
        "signature": "[class]android.widget.Button[resource_id]None[visible]True[text]Google Search[enabled,,]",
        "view_str": "7ca6e6231f59d98a1f6c1520b3110442",
        "bound_box": "42,372,168,493",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "6",
        "full_desc": "<button bound_box=42,372,168,493>Google Search</button>",
        "desc": "<button bound_box=42,372,168,493>Google Search</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            25
        ],
        "focused": false,
        "bounds": [
            [
                168,
                399
            ],
            [
                787,
                467
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 21,
        "temp_id": 24,
        "size": "619*68",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "49758e30796e16703a2ddfc5a8291621",
        "bound_box": "168,399,787,467",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": true,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                168,
                399
            ],
            [
                787,
                467
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "google",
        "class": "android.widget.EditText",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 24,
        "temp_id": 25,
        "size": "619*68",
        "signature": "[class]android.widget.EditText[resource_id]None[visible]True[text]google[enabled,,]",
        "view_str": "c66a0cb8395d2000a3aec7123b2b3c0a",
        "bound_box": "168,399,787,467",
        "content_free_signature": "[class]android.widget.EditText[resource_id]None[visible]True",
        "allowed_actions": [
            "touch",
            "set_text"
        ],
        "status": [],
        "local_id": "7",
        "full_desc": "<input bound_box=168,399,787,467>google</input>",
        "desc": "<input bound_box=168,399,787,467>google</input>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                784,
                372
            ],
            [
                913,
                493
            ]
        ],
        "resource_id": "tsuid_2-0yZ-jtAcyGptQPofi-iA8_3",
        "checked": false,
        "text": "Clear Search",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 21,
        "temp_id": 26,
        "size": "129*121",
        "signature": "[class]android.widget.Button[resource_id]tsuid_2-0yZ-jtAcyGptQPofi-iA8_3[visible]True[text]Clear Search[enabled,,]",
        "view_str": "e10fb784dbc7e3fdc32b95d03af85c41",
        "bound_box": "784,372,913,493",
        "content_free_signature": "[class]android.widget.Button[resource_id]tsuid_2-0yZ-jtAcyGptQPofi-iA8_3[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "8",
        "full_desc": "<button bound_box=784,372,913,493>Clear Search</button>",
        "desc": "<button bound_box=784,372,913,493>Clear Search</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                913,
                372
            ],
            [
                1042,
                493
            ]
        ],
        "resource_id": "Q7Ulpb",
        "checked": false,
        "text": "Search by voice",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 21,
        "temp_id": 27,
        "size": "129*121",
        "signature": "[class]android.widget.Button[resource_id]Q7Ulpb[visible]True[text]Search by voice[enabled,,]",
        "view_str": "dcae42d5d54c957e509b2cbcf3df083d",
        "bound_box": "913,372,1042,493",
        "content_free_signature": "[class]android.widget.Button[resource_id]Q7Ulpb[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "9",
        "full_desc": "<button bound_box=913,372,1042,493>Search by voice</button>",
        "desc": "<button bound_box=913,372,1042,493>Search by voice</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                488
            ],
            [
                1042,
                504
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 21,
        "temp_id": 28,
        "size": "1000*16",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "319dc4c1fce8d2135fa87d7a336ce880",
        "bound_box": "42,488,1042,504",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                498
            ],
            [
                1042,
                498
            ]
        ],
        "resource_id": "tophf",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 21,
        "temp_id": 29,
        "size": "1000*0",
        "signature": "[class]android.view.View[resource_id]tophf[visible]False[text][enabled,,]",
        "view_str": "771d31bd78b9924ad605a17894e97401",
        "bound_box": "42,498,1042,498",
        "content_free_signature": "[class]android.view.View[resource_id]tophf[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                210
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "lb",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 11,
        "temp_id": 30,
        "size": "1084*2066",
        "signature": "[class]android.view.View[resource_id]lb[visible]True[text][enabled,,]",
        "view_str": "83cc711d042cef233f6c4f47f3f0ce4c",
        "bound_box": "0,210,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]lb[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            32
        ],
        "focused": false,
        "bounds": [
            [
                0,
                493
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "gsr",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 11,
        "temp_id": 31,
        "size": "1084*1783",
        "signature": "[class]android.view.View[resource_id]gsr[visible]True[text][enabled,,]",
        "view_str": "44507fa9850f899a4a88ceef1007ea6e",
        "bound_box": "0,493,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]gsr[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            33
        ],
        "focused": false,
        "bounds": [
            [
                0,
                493
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "main",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 31,
        "temp_id": 32,
        "size": "1084*1783",
        "signature": "[class]android.view.View[resource_id]main[visible]True[text][enabled,,]",
        "view_str": "8bc3952a609d1b428b2d612a80cf8479",
        "bound_box": "0,493,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]main[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 12,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            36,
            93,
            96,
            627,
            631,
            635
        ],
        "focused": false,
        "bounds": [
            [
                0,
                493
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "cnt",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 32,
        "temp_id": 33,
        "size": "1084*1783",
        "signature": "[class]android.view.View[resource_id]cnt[visible]True[text][enabled,,]",
        "view_str": "4a7013c559ad7a0c15c624c8b6070fee",
        "bound_box": "0,493,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]cnt[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            35
        ],
        "focused": false,
        "bounds": [
            [
                0,
                779
            ],
            [
                1084,
                779
            ]
        ],
        "resource_id": "before-appbar",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 33,
        "temp_id": 34,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]before-appbar[visible]False[text][enabled,,]",
        "view_str": "b3805b05d67a83e46233fc15f98c31d6",
        "bound_box": "0,779,1084,779",
        "content_free_signature": "[class]android.view.View[resource_id]before-appbar[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                493
            ],
            [
                1084,
                493
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_14",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 34,
        "temp_id": 35,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_14[visible]False[text][enabled,,]",
        "view_str": "c8e7bafdf84b2315e79259535a0cde7a",
        "bound_box": "0,493,1084,493",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_14[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            37
        ],
        "focused": false,
        "bounds": [
            [
                0,
                493
            ],
            [
                1084,
                616
            ]
        ],
        "resource_id": "appbar",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 33,
        "temp_id": 36,
        "size": "1084*123",
        "signature": "[class]android.view.View[resource_id]appbar[visible]True[text][enabled,,]",
        "view_str": "b3df3162ead1deb32cfce687108ea66e",
        "bound_box": "0,493,1084,616",
        "content_free_signature": "[class]android.view.View[resource_id]appbar[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            38
        ],
        "focused": false,
        "bounds": [
            [
                0,
                493
            ],
            [
                1084,
                616
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Filters and Topics",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 36,
        "temp_id": 37,
        "size": "1084*123",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]Filters and Topics[enabled,,]",
        "view_str": "f58949e5596c90199cb7b11fea19361d",
        "bound_box": "0,493,1084,616",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "10",
        "full_desc": "<button bound_box=0,493,1084,616>Filters and Topics</button>",
        "desc": "<button bound_box=0,493,1084,616>Filters and Topics</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            39
        ],
        "focused": false,
        "bounds": [
            [
                0,
                493
            ],
            [
                1084,
                616
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 37,
        "temp_id": 38,
        "size": "1084*123",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "840617ff1a50d375e7286a04f1035a36",
        "bound_box": "0,493,1084,616",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            40
        ],
        "focused": false,
        "bounds": [
            [
                0,
                493
            ],
            [
                1084,
                616
            ]
        ],
        "resource_id": "bqHHPb",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 38,
        "temp_id": 39,
        "size": "1084*123",
        "signature": "[class]android.view.View[resource_id]bqHHPb[visible]True[text][enabled,,]",
        "view_str": "9f3baff1570d5ee8587e546ea85c4d31",
        "bound_box": "0,493,1084,616",
        "content_free_signature": "[class]android.view.View[resource_id]bqHHPb[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            41,
            42
        ],
        "focused": false,
        "bounds": [
            [
                0,
                493
            ],
            [
                1084,
                616
            ]
        ],
        "resource_id": "hdtb-sc",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 39,
        "temp_id": 40,
        "size": "1084*123",
        "signature": "[class]android.view.View[resource_id]hdtb-sc[visible]True[text][enabled,,]",
        "view_str": "0bc99b901e37df568a35d0f2964fdd72",
        "bound_box": "0,493,1084,616",
        "content_free_signature": "[class]android.view.View[resource_id]hdtb-sc[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "11",
        "full_desc": "<button bound_box=0,493,1084,616></button>",
        "desc": "<button bound_box=0,493,1084,616></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                504
            ],
            [
                5,
                509
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_26",
        "checked": false,
        "text": "Filters and Topics",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 40,
        "temp_id": 41,
        "size": "5*5",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_26[visible]True[text]Filters and Topics[enabled,,]",
        "view_str": "1be5f09c4e63d010573a2e5ee47e7766",
        "bound_box": "0,504,5,509",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_26[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "12",
        "full_desc": "<button bound_box=0,504,5,509>Filters and Topics</button>",
        "desc": "<button bound_box=0,504,5,509>Filters and Topics</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            43,
            44
        ],
        "focused": false,
        "bounds": [
            [
                0,
                504
            ],
            [
                1084,
                606
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 40,
        "temp_id": 42,
        "size": "1084*102",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "bcae97e111b0a1f26688f20c1b546c0a",
        "bound_box": "0,504,1084,606",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1018,
                504
            ],
            [
                1084,
                619
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 42,
        "temp_id": 43,
        "size": "66*115",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "5a936f9c11e73ada87403cc975278bbe",
        "bound_box": "1018,504,1084,619",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            45
        ],
        "focused": false,
        "bounds": [
            [
                0,
                504
            ],
            [
                1084,
                606
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 42,
        "temp_id": 44,
        "size": "1084*102",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "81b01df5e8113c75d102b2ed37651b90",
        "bound_box": "0,504,1084,606",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            46
        ],
        "focused": false,
        "bounds": [
            [
                0,
                504
            ],
            [
                1084,
                606
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": true,
        "selected": false,
        "long_clickable": false,
        "parent": 44,
        "temp_id": 45,
        "size": "1084*102",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "d553458087a577a50d3cb7d811e23440",
        "bound_box": "0,504,1084,606",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "scroll up",
            "scroll down",
            "scroll left",
            "scroll right"
        ],
        "status": [],
        "local_id": "13",
        "full_desc": "<button bound_box=0,504,1084,606></button>",
        "desc": "<button bound_box=0,504,1084,606></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            47
        ],
        "focused": false,
        "bounds": [
            [
                7,
                504
            ],
            [
                2488,
                606
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 45,
        "temp_id": 46,
        "size": "2481*102",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "9a6a2db084aa457b6a48b799d2a301be",
        "bound_box": "7,504,2488,606",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "14",
        "full_desc": "<button bound_box=7,504,2488,606></button>",
        "desc": "<button bound_box=7,504,2488,606></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [
            48
        ],
        "focused": false,
        "bounds": [
            [
                7,
                504
            ],
            [
                2488,
                606
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "All Images Videos News Short videos Forums Web Maps Books Flights Finance Search tools Feedback",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 46,
        "temp_id": 47,
        "size": "2481*102",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "31813636a686d21675dec202468f3435",
        "bound_box": "7,504,2488,606",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "15",
        "full_desc": "<button bound_box=7,504,2488,606>All Images Videos News Short videos Forums Web Map</button>",
        "desc": "<button bound_box=7,504,2488,606>All Images Videos News Short videos Forums Web Map</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 11,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            49,
            52,
            55,
            58,
            61,
            64,
            71,
            79
        ],
        "focused": false,
        "bounds": [
            [
                7,
                504
            ],
            [
                1913,
                606
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.widget.ListView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 47,
        "temp_id": 48,
        "size": "1906*102",
        "signature": "[class]android.widget.ListView[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "7f62770720a24c95c5332a7d0f2bacf6",
        "bound_box": "7,504,1913,606",
        "content_free_signature": "[class]android.widget.ListView[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            50
        ],
        "focused": false,
        "bounds": [
            [
                7,
                504
            ],
            [
                118,
                606
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 48,
        "temp_id": 49,
        "size": "111*102",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "95acf4b8430eb08b7a8a3f921ba76cd5",
        "bound_box": "7,504,118,606",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "16",
        "full_desc": "<button bound_box=7,504,118,606></button>",
        "desc": "<button bound_box=7,504,118,606></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": false,
        "content_description": "All, current page",
        "children": [
            51
        ],
        "focused": false,
        "bounds": [
            [
                7,
                504
            ],
            [
                118,
                606
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "All",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 49,
        "temp_id": 50,
        "size": "111*102",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]All[,,]",
        "view_str": "766f37981b3cdd08673817c9ce5838f4",
        "bound_box": "7,504,118,606",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "17",
        "full_desc": "<button alt='All, current page' bound_box=7,504,118,606>All</button>",
        "desc": "<button alt='All, current page' bound_box=7,504,118,606>All</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                532
            ],
            [
                86,
                580
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "All",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 50,
        "temp_id": 51,
        "size": "44*48",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]True[text]All[enabled,,]",
        "view_str": "5d465b676cb1050909fc6f331e7622e7",
        "bound_box": "42,532,86,580",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "18",
        "full_desc": "<button bound_box=42,532,86,580>All</button>",
        "desc": "<button bound_box=42,532,86,580>All</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            53
        ],
        "focused": false,
        "bounds": [
            [
                115,
                504
            ],
            [
                304,
                606
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 48,
        "temp_id": 52,
        "size": "189*102",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "9e57af87052be3077496b0d5fe6b3a8c",
        "bound_box": "115,504,304,606",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "19",
        "full_desc": "<button bound_box=115,504,304,606></button>",
        "desc": "<button bound_box=115,504,304,606></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Images",
        "children": [
            54
        ],
        "focused": false,
        "bounds": [
            [
                115,
                504
            ],
            [
                304,
                598
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 52,
        "temp_id": 53,
        "size": "189*94",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "e8fcc4c48c10a3aadeba2b7a18ae5588",
        "bound_box": "115,504,304,598",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "20",
        "full_desc": "<button alt='Images' bound_box=115,504,304,598></button>",
        "desc": "<button alt='Images' bound_box=115,504,304,598></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                147,
                532
            ],
            [
                270,
                580
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Images",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 53,
        "temp_id": 54,
        "size": "123*48",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]True[text]Images[enabled,,]",
        "view_str": "6f733433a1f6f5c82b3b418f51c02242",
        "bound_box": "147,532,270,580",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "21",
        "full_desc": "<button bound_box=147,532,270,580>Images</button>",
        "desc": "<button bound_box=147,532,270,580>Images</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            56
        ],
        "focused": false,
        "bounds": [
            [
                299,
                504
            ],
            [
                480,
                606
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 48,
        "temp_id": 55,
        "size": "181*102",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "9e57af87052be3077496b0d5fe6b3a8c",
        "bound_box": "299,504,480,606",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "22",
        "full_desc": "<button bound_box=299,504,480,606></button>",
        "desc": "<button bound_box=299,504,480,606></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Videos",
        "children": [
            57
        ],
        "focused": false,
        "bounds": [
            [
                299,
                504
            ],
            [
                480,
                598
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 55,
        "temp_id": 56,
        "size": "181*94",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "bfde6871e1c8e01857c0b3879bf5507e",
        "bound_box": "299,504,480,598",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "23",
        "full_desc": "<button alt='Videos' bound_box=299,504,480,598></button>",
        "desc": "<button alt='Videos' bound_box=299,504,480,598></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                330,
                532
            ],
            [
                448,
                580
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Videos",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 56,
        "temp_id": 57,
        "size": "118*48",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]True[text]Videos[enabled,,]",
        "view_str": "165ef3e8008945d87fafc1ecf5ce6c0e",
        "bound_box": "330,532,448,580",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "24",
        "full_desc": "<button bound_box=330,532,448,580>Videos</button>",
        "desc": "<button bound_box=330,532,448,580>Videos</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            59
        ],
        "focused": false,
        "bounds": [
            [
                475,
                504
            ],
            [
                635,
                606
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 48,
        "temp_id": 58,
        "size": "160*102",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "9e57af87052be3077496b0d5fe6b3a8c",
        "bound_box": "475,504,635,606",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "25",
        "full_desc": "<button bound_box=475,504,635,606></button>",
        "desc": "<button bound_box=475,504,635,606></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "News",
        "children": [
            60
        ],
        "focused": false,
        "bounds": [
            [
                475,
                504
            ],
            [
                635,
                598
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 58,
        "temp_id": 59,
        "size": "160*94",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "1a3d2b070be5b48d5fb405fc9aaa2c5a",
        "bound_box": "475,504,635,598",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "26",
        "full_desc": "<button alt='News' bound_box=475,504,635,598></button>",
        "desc": "<button alt='News' bound_box=475,504,635,598></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                506,
                532
            ],
            [
                601,
                580
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "News",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 59,
        "temp_id": 60,
        "size": "95*48",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]True[text]News[enabled,,]",
        "view_str": "4ce1b477295beea63532ed8be1c66550",
        "bound_box": "506,532,601,580",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "27",
        "full_desc": "<button bound_box=506,532,601,580>News</button>",
        "desc": "<button bound_box=506,532,601,580>News</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            62
        ],
        "focused": false,
        "bounds": [
            [
                630,
                504
            ],
            [
                903,
                606
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 48,
        "temp_id": 61,
        "size": "273*102",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "9e57af87052be3077496b0d5fe6b3a8c",
        "bound_box": "630,504,903,606",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "28",
        "full_desc": "<button bound_box=630,504,903,606></button>",
        "desc": "<button bound_box=630,504,903,606></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Short videos",
        "children": [
            63
        ],
        "focused": false,
        "bounds": [
            [
                630,
                504
            ],
            [
                903,
                598
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 61,
        "temp_id": 62,
        "size": "273*94",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "231b92115651c82ce5fe0c97ff6a17c1",
        "bound_box": "630,504,903,598",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "29",
        "full_desc": "<button alt='Short videos' bound_box=630,504,903,598></button>",
        "desc": "<button alt='Short videos' bound_box=630,504,903,598></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                661,
                532
            ],
            [
                871,
                580
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Short videos",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 62,
        "temp_id": 63,
        "size": "210*48",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]True[text]Short videos[enabled,,]",
        "view_str": "86d7ef1fc0b56fa42cd5f5109e7ff820",
        "bound_box": "661,532,871,580",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "30",
        "full_desc": "<button bound_box=661,532,871,580>Short videos</button>",
        "desc": "<button bound_box=661,532,871,580>Short videos</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            65
        ],
        "focused": false,
        "bounds": [
            [
                900,
                504
            ],
            [
                1092,
                606
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 48,
        "temp_id": 64,
        "size": "192*102",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "9e57af87052be3077496b0d5fe6b3a8c",
        "bound_box": "900,504,1092,606",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "31",
        "full_desc": "<button bound_box=900,504,1092,606></button>",
        "desc": "<button bound_box=900,504,1092,606></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Forums",
        "children": [
            66
        ],
        "focused": false,
        "bounds": [
            [
                900,
                504
            ],
            [
                1092,
                598
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 64,
        "temp_id": 65,
        "size": "192*94",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "de6e97461cc634e15ead10a340a02abe",
        "bound_box": "900,504,1092,598",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "32",
        "full_desc": "<button alt='Forums' bound_box=900,504,1092,598></button>",
        "desc": "<button alt='Forums' bound_box=900,504,1092,598></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                931,
                532
            ],
            [
                1060,
                580
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Forums",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 65,
        "temp_id": 66,
        "size": "129*48",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]True[text]Forums[enabled,,]",
        "view_str": "86e2d8b35ab4ebb4f0c5bb8f76368d80",
        "bound_box": "931,532,1060,580",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "33",
        "full_desc": "<button bound_box=931,532,1060,580>Forums</button>",
        "desc": "<button bound_box=931,532,1060,580>Forums</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            68
        ],
        "focused": false,
        "bounds": [
            [
                1089,
                504
            ],
            [
                1228,
                606
            ]
        ],
        "resource_id": "2-0yZ-jtAcyGptQPofi-iA8__14",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 48,
        "temp_id": 67,
        "size": "139*102",
        "signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__14[visible]False[text][enabled,,]",
        "view_str": "f06c29e821a3f708551d120b0d3077d7",
        "bound_box": "1089,504,1228,606",
        "content_free_signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__14[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            69
        ],
        "focused": false,
        "bounds": [
            [
                1089,
                504
            ],
            [
                1228,
                606
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 67,
        "temp_id": 68,
        "size": "139*102",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "c76e1f7dca5785a80340497df0fabc04",
        "bound_box": "1089,504,1228,606",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Web",
        "children": [
            70
        ],
        "focused": false,
        "bounds": [
            [
                1089,
                504
            ],
            [
                1228,
                598
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 68,
        "temp_id": 69,
        "size": "139*94",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "5db444333d83583a2cd69cd32b5fa7aa",
        "bound_box": "1089,504,1228,598",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1120,
                532
            ],
            [
                1194,
                580
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Web",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 69,
        "temp_id": 70,
        "size": "74*48",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]Web[enabled,,]",
        "view_str": "a631fc5ffa1086f18092db3605042ff0",
        "bound_box": "1120,532,1194,580",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            72
        ],
        "focused": false,
        "bounds": [
            [
                1223,
                504
            ],
            [
                1380,
                606
            ]
        ],
        "resource_id": "2-0yZ-jtAcyGptQPofi-iA8__15",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 48,
        "temp_id": 71,
        "size": "157*102",
        "signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__15[visible]False[text][enabled,,]",
        "view_str": "2f4bc86c82acbd5545ede56ac7d6eea0",
        "bound_box": "1223,504,1380,606",
        "content_free_signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__15[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            73
        ],
        "focused": false,
        "bounds": [
            [
                1223,
                504
            ],
            [
                1380,
                606
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 71,
        "temp_id": 72,
        "size": "157*102",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "529c25757adbb96bd38f69b478e3f8df",
        "bound_box": "1223,504,1380,606",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Maps",
        "children": [
            74
        ],
        "focused": false,
        "bounds": [
            [
                1223,
                504
            ],
            [
                1380,
                598
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 72,
        "temp_id": 73,
        "size": "157*94",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "a03ca3d5c550fe6e10e5054a02d7c441",
        "bound_box": "1223,504,1380,598",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1254,
                532
            ],
            [
                1349,
                580
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Maps",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 73,
        "temp_id": 74,
        "size": "95*48",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]Maps[enabled,,]",
        "view_str": "21b350e96d18de4b59fa4198b0aa1a48",
        "bound_box": "1254,532,1349,580",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            76
        ],
        "focused": false,
        "bounds": [
            [
                1378,
                504
            ],
            [
                1546,
                606
            ]
        ],
        "resource_id": "2-0yZ-jtAcyGptQPofi-iA8__16",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 48,
        "temp_id": 75,
        "size": "168*102",
        "signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__16[visible]False[text][enabled,,]",
        "view_str": "88c695709f39c1cbc38982193976fc25",
        "bound_box": "1378,504,1546,606",
        "content_free_signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__16[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            77
        ],
        "focused": false,
        "bounds": [
            [
                1378,
                504
            ],
            [
                1546,
                606
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 75,
        "temp_id": 76,
        "size": "168*102",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "86c6a412d73af8fd44ffe93e433ba16b",
        "bound_box": "1378,504,1546,606",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Books",
        "children": [
            78
        ],
        "focused": false,
        "bounds": [
            [
                1378,
                504
            ],
            [
                1546,
                598
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 76,
        "temp_id": 77,
        "size": "168*94",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "9b9a823005b27e461b2839af84c59491",
        "bound_box": "1378,504,1546,598",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1409,
                532
            ],
            [
                1517,
                580
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Books",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 77,
        "temp_id": 78,
        "size": "108*48",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]Books[enabled,,]",
        "view_str": "9bae2665c7f7e6fa896bbaf339cda447",
        "bound_box": "1409,532,1517,580",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            80
        ],
        "focused": false,
        "bounds": [
            [
                1543,
                504
            ],
            [
                1722,
                606
            ]
        ],
        "resource_id": "2-0yZ-jtAcyGptQPofi-iA8__17",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 48,
        "temp_id": 79,
        "size": "179*102",
        "signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__17[visible]False[text][enabled,,]",
        "view_str": "85f87e456a854e72f0bfd3925f5921ea",
        "bound_box": "1543,504,1722,606",
        "content_free_signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__17[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            81
        ],
        "focused": false,
        "bounds": [
            [
                1543,
                504
            ],
            [
                1722,
                606
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 79,
        "temp_id": 80,
        "size": "179*102",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "acf249182b99ce5d3ee8478fedd5f4eb",
        "bound_box": "1543,504,1722,606",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Flights",
        "children": [
            82
        ],
        "focused": false,
        "bounds": [
            [
                1543,
                504
            ],
            [
                1722,
                598
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 80,
        "temp_id": 81,
        "size": "179*94",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "eb36d6585906ad36fd5c1c2ac387245b",
        "bound_box": "1543,504,1722,598",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1575,
                532
            ],
            [
                1690,
                580
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Flights",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 81,
        "temp_id": 82,
        "size": "115*48",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]Flights[enabled,,]",
        "view_str": "55a6aa2810c4a09af135ddb03436a776",
        "bound_box": "1575,532,1690,580",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            84
        ],
        "focused": false,
        "bounds": [
            [
                1719,
                504
            ],
            [
                1913,
                606
            ]
        ],
        "resource_id": "2-0yZ-jtAcyGptQPofi-iA8__19",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 48,
        "temp_id": 83,
        "size": "194*102",
        "signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__19[visible]False[text][enabled,,]",
        "view_str": "6844eed566f1a6da4af571c5df687381",
        "bound_box": "1719,504,1913,606",
        "content_free_signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__19[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            85
        ],
        "focused": false,
        "bounds": [
            [
                1719,
                504
            ],
            [
                1913,
                606
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 83,
        "temp_id": 84,
        "size": "194*102",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "5034b6764f4a4224313e47e0c76ae04b",
        "bound_box": "1719,504,1913,606",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Finance",
        "children": [
            86
        ],
        "focused": false,
        "bounds": [
            [
                1719,
                504
            ],
            [
                1913,
                598
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 84,
        "temp_id": 85,
        "size": "194*94",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "7494c8cbf1f44e09f670b6aa448ca814",
        "bound_box": "1719,504,1913,598",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1750,
                532
            ],
            [
                1882,
                580
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Finance",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 85,
        "temp_id": 86,
        "size": "132*48",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]Finance[enabled,,]",
        "view_str": "f8c9706fc424d0269a9e90b24583f4e8",
        "bound_box": "1750,532,1882,580",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            88
        ],
        "focused": false,
        "bounds": [
            [
                1911,
                519
            ],
            [
                2488,
                593
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.widget.ListView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 47,
        "temp_id": 87,
        "size": "577*74",
        "signature": "[class]android.widget.ListView[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "a491d2b91b3243f6489fb46b0ca1e023",
        "bound_box": "1911,519,2488,593",
        "content_free_signature": "[class]android.widget.ListView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            89,
            90
        ],
        "focused": false,
        "bounds": [
            [
                1921,
                525
            ],
            [
                2462,
                593
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_29",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 87,
        "temp_id": 88,
        "size": "541*68",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_29[visible]False[text][enabled,,]",
        "view_str": "84a77efe9c03ac1990e84da94d205b5d",
        "bound_box": "1921,525,2462,593",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_29[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1924,
                525
            ],
            [
                2215,
                593
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Search tools",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 88,
        "temp_id": 89,
        "size": "291*68",
        "signature": "[class]android.widget.Button[resource_id]None[visible]False[text]Search tools[enabled,,]",
        "view_str": "a47089b9ce963b3798a5da64274ad595",
        "bound_box": "1924,525,2215,593",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Feedback",
        "children": [
            91
        ],
        "focused": false,
        "bounds": [
            [
                2215,
                525
            ],
            [
                2462,
                593
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 88,
        "temp_id": 90,
        "size": "247*68",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "327014e334daf3c245d135e747380531",
        "bound_box": "2215,525,2462,593",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                2257,
                535
            ],
            [
                2420,
                580
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Feedback",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 90,
        "temp_id": 91,
        "size": "163*45",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]Feedback[enabled,,]",
        "view_str": "7c093b8ddc7604d041dc25b3152c56bf",
        "bound_box": "2257,535,2420,580",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                900
            ],
            [
                1084,
                900
            ]
        ],
        "resource_id": "easter-egg",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 33,
        "temp_id": 92,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]easter-egg[visible]False[text][enabled,,]",
        "view_str": "cec494d7be349d897aab8068d7988436",
        "bound_box": "0,900,1084,900",
        "content_free_signature": "[class]android.view.View[resource_id]easter-egg[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                614
            ],
            [
                1084,
                614
            ]
        ],
        "resource_id": "appbar-previews",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 33,
        "temp_id": 93,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]appbar-previews[visible]False[text][enabled,,]",
        "view_str": "9b967e9ddd375c0bb52a0057d9a641a6",
        "bound_box": "0,614,1084,614",
        "content_free_signature": "[class]android.view.View[resource_id]appbar-previews[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            95
        ],
        "focused": false,
        "bounds": [
            [
                0,
                900
            ],
            [
                1084,
                900
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_34",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 33,
        "temp_id": 94,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_34[visible]False[text][enabled,,]",
        "view_str": "8434a82fda1d13630c75c37041003368",
        "bound_box": "0,900,1084,900",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_34[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                614
            ],
            [
                1084,
                614
            ]
        ],
        "resource_id": "arc-stev",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 94,
        "temp_id": 95,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]arc-stev[visible]False[text][enabled,,]",
        "view_str": "4241bc42aa2d7d5fa442af7e7bc83f97",
        "bound_box": "0,614,1084,614",
        "content_free_signature": "[class]android.view.View[resource_id]arc-stev[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 6,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            100,
            101,
            578
        ],
        "focused": false,
        "bounds": [
            [
                0,
                614
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "center_col",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 33,
        "temp_id": 96,
        "size": "1084*1662",
        "signature": "[class]android.view.View[resource_id]center_col[visible]True[text][enabled,,]",
        "view_str": "cbc7ff36a479078ba0b4943e240123b8",
        "bound_box": "0,614,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]center_col[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            98
        ],
        "focused": false,
        "bounds": [
            [
                0,
                900
            ],
            [
                1084,
                900
            ]
        ],
        "resource_id": "taw",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 96,
        "temp_id": 97,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]taw[visible]False[text][enabled,,]",
        "view_str": "9abd3ed73d87fc9a539155f53413ed4d",
        "bound_box": "0,900,1084,900",
        "content_free_signature": "[class]android.view.View[resource_id]taw[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            99
        ],
        "focused": false,
        "bounds": [
            [
                0,
                900
            ],
            [
                1084,
                900
            ]
        ],
        "resource_id": "tvcap",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 97,
        "temp_id": 98,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]tvcap[visible]False[text][enabled,,]",
        "view_str": "de0b05bc033a5c0a733db5126bb600b7",
        "bound_box": "0,900,1084,900",
        "content_free_signature": "[class]android.view.View[resource_id]tvcap[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                900
            ],
            [
                1084,
                900
            ]
        ],
        "resource_id": "tads",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 98,
        "temp_id": 99,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]tads[visible]False[text][enabled,,]",
        "view_str": "efd9201f0149de5c2148918eebb8faf2",
        "bound_box": "0,900,1084,900",
        "content_free_signature": "[class]android.view.View[resource_id]tads[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                614
            ],
            [
                1084,
                614
            ]
        ],
        "resource_id": "topstuff",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 96,
        "temp_id": 100,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]topstuff[visible]False[text][enabled,,]",
        "view_str": "42184fd2255ae532270775a3e8404c13",
        "bound_box": "0,614,1084,614",
        "content_free_signature": "[class]android.view.View[resource_id]topstuff[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            102,
            103
        ],
        "focused": false,
        "bounds": [
            [
                0,
                614
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 96,
        "temp_id": 101,
        "size": "1084*1662",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "ace6b34843a4bae5836ecbabe3bd066b",
        "bound_box": "0,614,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "34",
        "full_desc": "<button bound_box=0,614,1084,2276></button>",
        "desc": "<button bound_box=0,614,1084,2276></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                614
            ],
            [
                5,
                619
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Search Results",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 101,
        "temp_id": 102,
        "size": "5*5",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]Search Results[enabled,,]",
        "view_str": "69200426579bcbd0bcdbafd56018361f",
        "bound_box": "0,614,5,619",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "35",
        "full_desc": "<button bound_box=0,614,5,619>Search Results</button>",
        "desc": "<button bound_box=0,614,5,619>Search Results</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 13,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            104,
            236,
            237,
            294,
            397,
            413,
            513
        ],
        "focused": false,
        "bounds": [
            [
                0,
                614
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "rso",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 101,
        "temp_id": 103,
        "size": "1084*1662",
        "signature": "[class]android.view.View[resource_id]rso[visible]True[text][enabled,,]",
        "view_str": "ca0a84a31951a6e816465a5076c7de84",
        "bound_box": "0,614,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]rso[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            107
        ],
        "focused": false,
        "bounds": [
            [
                0,
                614
            ],
            [
                1084,
                2218
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 103,
        "temp_id": 104,
        "size": "1084*1604",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "74eeb3cb7e20bac9e3829ab6d64179d2",
        "bound_box": "0,614,1084,2218",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "36",
        "full_desc": "<button bound_box=0,614,1084,2218></button>",
        "desc": "<button bound_box=0,614,1084,2218></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            106
        ],
        "focused": false,
        "bounds": [
            [
                0,
                900
            ],
            [
                1084,
                900
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_41",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 104,
        "temp_id": 105,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_41[visible]False[text][enabled,,]",
        "view_str": "37d45efae8e853bcbcb9660350fb18e3",
        "bound_box": "0,900,1084,900",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_41[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                614
            ],
            [
                1084,
                614
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_44",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 105,
        "temp_id": 106,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_44[visible]False[text][enabled,,]",
        "view_str": "c25f2c6ebf6c151de7947a4544b5bd38",
        "bound_box": "0,614,1084,614",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_44[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            108,
            119
        ],
        "focused": false,
        "bounds": [
            [
                0,
                614
            ],
            [
                1084,
                2218
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_33",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 104,
        "temp_id": 107,
        "size": "1084*1604",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_33[visible]True[text][enabled,,]",
        "view_str": "ddafb2b7603a5fe8ed58cd4ffbaf98c5",
        "bound_box": "0,614,1084,2218",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_33[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            109
        ],
        "focused": false,
        "bounds": [
            [
                0,
                614
            ],
            [
                1084,
                847
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 107,
        "temp_id": 108,
        "size": "1084*233",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "5fdb5e75c81352787920422d344e2236",
        "bound_box": "0,614,1084,847",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "37",
        "full_desc": "<button bound_box=0,614,1084,847></button>",
        "desc": "<button bound_box=0,614,1084,847></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            110
        ],
        "focused": false,
        "bounds": [
            [
                0,
                614
            ],
            [
                1084,
                847
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 108,
        "temp_id": 109,
        "size": "1084*233",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "0d2f016c542ab4080f85faac3b816a3d",
        "bound_box": "0,614,1084,847",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 4,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            111,
            112,
            113,
            118
        ],
        "focused": false,
        "bounds": [
            [
                42,
                656
            ],
            [
                1042,
                826
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 109,
        "temp_id": 110,
        "size": "1000*170",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "05940aabb17f4ea12911706ef595e3b8",
        "bound_box": "42,656,1042,826",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                656
            ],
            [
                771,
                742
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 110,
        "temp_id": 111,
        "size": "729*86",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]Google[enabled,,]",
        "view_str": "a472a168d3d0b889159a312766b38489",
        "bound_box": "42,656,771,742",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "38",
        "full_desc": "<button bound_box=42,656,771,742>Google</button>",
        "desc": "<button bound_box=42,656,771,742>Google</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                750
            ],
            [
                845,
                805
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "IT corporation",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 110,
        "temp_id": 112,
        "size": "803*55",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]IT corporation[enabled,,]",
        "view_str": "ecaac994d225c18d54866bd1f7e5377a",
        "bound_box": "42,750,845,805",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "39",
        "full_desc": "<button bound_box=42,750,845,805>IT corporation</button>",
        "desc": "<button bound_box=42,750,845,805>IT corporation</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            114
        ],
        "focused": false,
        "bounds": [
            [
                745,
                679
            ],
            [
                845,
                766
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 110,
        "temp_id": 113,
        "size": "100*87",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "09b3f30676f9fdf106a30263d17d1bae",
        "bound_box": "745,679,845,766",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            115
        ],
        "focused": false,
        "bounds": [
            [
                766,
                666
            ],
            [
                871,
                753
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 113,
        "temp_id": 114,
        "size": "105*87",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "e530e321098b8351a93b37b6850463e6",
        "bound_box": "766,666,871,753",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            116
        ],
        "focused": false,
        "bounds": [
            [
                766,
                666
            ],
            [
                871,
                753
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 114,
        "temp_id": 115,
        "size": "105*87",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "685f2939beae32601b9f87b7377733c9",
        "bound_box": "766,666,871,753",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            117
        ],
        "focused": false,
        "bounds": [
            [
                766,
                666
            ],
            [
                871,
                753
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 115,
        "temp_id": 116,
        "size": "105*87",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "615e9e94219242a2da29369837581cde",
        "bound_box": "766,666,871,753",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                766,
                666
            ],
            [
                871,
                753
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "More options",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 116,
        "temp_id": 117,
        "size": "105*87",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]More options[enabled,,]",
        "view_str": "a141042b4988683dc5875c2a95ea16e0",
        "bound_box": "766,666,871,753",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "40",
        "full_desc": "<button bound_box=766,666,871,753>More options</button>",
        "desc": "<button bound_box=766,666,871,753>More options</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                871,
                656
            ],
            [
                1042,
                826
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Thumbnail image for Google",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 110,
        "temp_id": 118,
        "size": "171*170",
        "signature": "[class]android.widget.Button[resource_id]None[visible]True[text]Thumbnail image for Google[enabled,,]",
        "view_str": "c79824d3a8499f484c0d48be34b8c00c",
        "bound_box": "871,656,1042,826",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "41",
        "full_desc": "<button bound_box=871,656,1042,826>Thumbnail image for Google</button>",
        "desc": "<button bound_box=871,656,1042,826>Thumbnail image for Google</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            120,
            230
        ],
        "focused": false,
        "bounds": [
            [
                0,
                845
            ],
            [
                1084,
                2218
            ]
        ],
        "resource_id": "jobWhd",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 107,
        "temp_id": 119,
        "size": "1084*1373",
        "signature": "[class]android.view.View[resource_id]jobWhd[visible]True[text][enabled,,]",
        "view_str": "34f862cdf2ae94b0f2827bb56099bb2a",
        "bound_box": "0,845,1084,2218",
        "content_free_signature": "[class]android.view.View[resource_id]jobWhd[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            121,
            122
        ],
        "focused": false,
        "bounds": [
            [
                0,
                845
            ],
            [
                1084,
                2023
            ]
        ],
        "resource_id": "kp-wp-tab-cont-overview",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 119,
        "temp_id": 120,
        "size": "1084*1178",
        "signature": "[class]android.view.View[resource_id]kp-wp-tab-cont-overview[visible]True[text][enabled,,]",
        "view_str": "6693ba27acfbb8790d7a77631fc6c996",
        "bound_box": "0,845,1084,2023",
        "content_free_signature": "[class]android.view.View[resource_id]kp-wp-tab-cont-overview[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "42",
        "full_desc": "<button bound_box=0,845,1084,2023></button>",
        "desc": "<button bound_box=0,845,1084,2023></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                845
            ],
            [
                5,
                850
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Main Results",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 120,
        "temp_id": 121,
        "size": "5*5",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]Main Results[enabled,,]",
        "view_str": "f8688292307f023e5c256e1b44fb8866",
        "bound_box": "0,845,5,850",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "43",
        "full_desc": "<button bound_box=0,845,5,850>Main Results</button>",
        "desc": "<button bound_box=0,845,5,850>Main Results</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            123
        ],
        "focused": false,
        "bounds": [
            [
                0,
                845
            ],
            [
                1084,
                2023
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 120,
        "temp_id": 122,
        "size": "1084*1178",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "834107f1e27825fd383278f53a4478a6",
        "bound_box": "0,845,1084,2023",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 4,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            124,
            125,
            221,
            222
        ],
        "focused": false,
        "bounds": [
            [
                0,
                824
            ],
            [
                1084,
                2026
            ]
        ],
        "resource_id": "kp-wp-tab-overview",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 122,
        "temp_id": 123,
        "size": "1084*1202",
        "signature": "[class]android.view.View[resource_id]kp-wp-tab-overview[visible]True[text][enabled,,]",
        "view_str": "13a346aa1690f6711490ddc33782c846",
        "bound_box": "0,824,1084,2026",
        "content_free_signature": "[class]android.view.View[resource_id]kp-wp-tab-overview[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "44",
        "full_desc": "<button bound_box=0,824,1084,2026></button>",
        "desc": "<button bound_box=0,824,1084,2026></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                824
            ],
            [
                1084,
                2026
            ]
        ],
        "resource_id": "fld_2-0yZ-jtAcyGptQPofi-iA8_1",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 123,
        "temp_id": 124,
        "size": "1084*1202",
        "signature": "[class]android.view.View[resource_id]fld_2-0yZ-jtAcyGptQPofi-iA8_1[visible]True[text][enabled,,]",
        "view_str": "552cb2703000ead469b08da63efbf793",
        "bound_box": "0,824,1084,2026",
        "content_free_signature": "[class]android.view.View[resource_id]fld_2-0yZ-jtAcyGptQPofi-iA8_1[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 3,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            126,
            157,
            158
        ],
        "focused": false,
        "bounds": [
            [
                0,
                824
            ],
            [
                1084,
                1727
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 123,
        "temp_id": 125,
        "size": "1084*903",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "c2b94d04b001b7f070411041e251b2d1",
        "bound_box": "0,824,1084,1727",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "45",
        "full_desc": "<button bound_box=0,824,1084,1727></button>",
        "desc": "<button bound_box=0,824,1084,1727></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            127,
            137
        ],
        "focused": false,
        "bounds": [
            [
                0,
                824
            ],
            [
                1084,
                1454
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_48",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 125,
        "temp_id": 126,
        "size": "1084*630",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_48[visible]True[text][enabled,,]",
        "view_str": "48e677623d27fe4914aab2756d2945bf",
        "bound_box": "0,824,1084,1454",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_48[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            128
        ],
        "focused": false,
        "bounds": [
            [
                42,
                866
            ],
            [
                1042,
                1120
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 126,
        "temp_id": 127,
        "size": "1000*254",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "e76ccd97ceb7e3e5fb8082e3ba4dde28",
        "bound_box": "42,866,1042,1120",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            129
        ],
        "focused": false,
        "bounds": [
            [
                42,
                866
            ],
            [
                1042,
                1120
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 127,
        "temp_id": 128,
        "size": "1000*254",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "ac94a2d925c06296926fff54f0722688",
        "bound_box": "42,866,1042,1120",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            130
        ],
        "focused": false,
        "bounds": [
            [
                42,
                866
            ],
            [
                1042,
                1120
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 128,
        "temp_id": 129,
        "size": "1000*254",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "73665398e88c1370b28efd00eb02d22a",
        "bound_box": "42,866,1042,1120",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "46",
        "full_desc": "<button bound_box=42,866,1042,1120></button>",
        "desc": "<button bound_box=42,866,1042,1120></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [
            131,
            135
        ],
        "focused": false,
        "bounds": [
            [
                55,
                882
            ],
            [
                1026,
                1105
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google LLC is an American-based multinational corporation and technology company focusing on online advertising, search engine technology, cloud computing, computer software, quantum computing, e-commerce, consumer electronics, and artificial intelligence.Wikipedia",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 129,
        "temp_id": 130,
        "size": "971*223",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "a65731cd6f77165c14976ea13893ec75",
        "bound_box": "55,882,1026,1105",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "47",
        "full_desc": "<button bound_box=55,882,1026,1105>Google LLC is an American-based multinational corp</button>",
        "desc": "<button bound_box=55,882,1026,1105>Google LLC is an American-based multinational corp</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            132,
            133
        ],
        "focused": false,
        "bounds": [
            [
                70,
                897
            ],
            [
                947,
                1089
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 130,
        "temp_id": 131,
        "size": "877*192",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "077c0f7cc3dad99eb9aaa889ca2efa48",
        "bound_box": "70,897,947,1089",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                70,
                897
            ],
            [
                945,
                1183
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google LLC is an American-based multinational corporation and technology company focusing on online advertising, search engine technology, cloud computing, computer software, quantum computing, e-commerce, consumer electronics, and artificial intelligence.",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 131,
        "temp_id": 132,
        "size": "875*286",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "f405ac51f91f58d70a5a80251b7c3145",
        "bound_box": "70,897,945,1183",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "48",
        "full_desc": "<button bound_box=70,897,945,1183>Google LLC is an American-based multinational corp</button>",
        "desc": "<button bound_box=70,897,945,1183>Google LLC is an American-based multinational corp</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Wikipedia",
        "children": [
            134
        ],
        "focused": false,
        "bounds": [
            [
                727,
                1039
            ],
            [
                947,
                1089
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 131,
        "temp_id": 133,
        "size": "220*50",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "193984b3881509f8f1519434e4c26e88",
        "bound_box": "727,1039,947,1089",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "49",
        "full_desc": "<button alt='Wikipedia' bound_box=727,1039,947,1089></button>",
        "desc": "<button alt='Wikipedia' bound_box=727,1039,947,1089></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                727,
                1039
            ],
            [
                947,
                1089
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Wikipedia",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 133,
        "temp_id": 134,
        "size": "220*50",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]Wikipedia[enabled,,]",
        "view_str": "b67056e604722817b9154736f70e365b",
        "bound_box": "727,1039,947,1089",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "50",
        "full_desc": "<button bound_box=727,1039,947,1089>Wikipedia</button>",
        "desc": "<button bound_box=727,1039,947,1089>Wikipedia</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            136
        ],
        "focused": false,
        "bounds": [
            [
                884,
                824
            ],
            [
                1078,
                1026
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 130,
        "temp_id": 135,
        "size": "194*202",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "0fa85247464063f700215b52bb931df2",
        "bound_box": "884,824,1078,1026",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                947,
                887
            ],
            [
                1015,
                952
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.widget.Image",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 135,
        "temp_id": 136,
        "size": "68*65",
        "signature": "[class]android.widget.Image[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "ac2fdfa80310c99a6e1153c8f8910d51",
        "bound_box": "947,887,1015,952",
        "content_free_signature": "[class]android.widget.Image[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            138,
            146
        ],
        "focused": false,
        "bounds": [
            [
                42,
                1149
            ],
            [
                1042,
                1412
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 126,
        "temp_id": 137,
        "size": "1000*263",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "bdb1552f164426f19bca7d65f0abc8df",
        "bound_box": "42,1149,1042,1412",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            139
        ],
        "focused": false,
        "bounds": [
            [
                42,
                1149
            ],
            [
                527,
                1412
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 137,
        "temp_id": 138,
        "size": "485*263",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "ac94a2d925c06296926fff54f0722688",
        "bound_box": "42,1149,527,1412",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            140
        ],
        "focused": false,
        "bounds": [
            [
                42,
                1149
            ],
            [
                527,
                1412
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 138,
        "temp_id": 139,
        "size": "485*263",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "73665398e88c1370b28efd00eb02d22a",
        "bound_box": "42,1149,527,1412",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "51",
        "full_desc": "<button bound_box=42,1149,527,1412></button>",
        "desc": "<button bound_box=42,1149,527,1412></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Age 26 years September 4, 1998",
        "children": [
            141
        ],
        "focused": false,
        "bounds": [
            [
                42,
                1149
            ],
            [
                527,
                1412
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 139,
        "temp_id": 140,
        "size": "485*263",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "e95d52f3c46d74e24fc4d2ac0a0bc582",
        "bound_box": "42,1149,527,1412",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "52",
        "full_desc": "<button alt='Age 26 years September 4, 1998' bound_box=42,1149,527,1412></button>",
        "desc": "<button alt='Age 26 years September 4, 1998' bound_box=42,1149,527,1412></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            142,
            143
        ],
        "focused": false,
        "bounds": [
            [
                42,
                1149
            ],
            [
                527,
                1412
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 140,
        "temp_id": 141,
        "size": "485*263",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "60a6bd8739bf4a61f375a0a6d05ffb04",
        "bound_box": "42,1149,527,1412",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                70,
                1178
            ],
            [
                496,
                1257
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_51",
        "checked": false,
        "text": "Age",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 141,
        "temp_id": 142,
        "size": "426*79",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_51[visible]True[text]Age[enabled,,]",
        "view_str": "c5bf79a7724ee7f93fae24bc8b14a170",
        "bound_box": "70,1178,496,1257",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_51[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "53",
        "full_desc": "<button bound_box=70,1178,496,1257>Age</button>",
        "desc": "<button bound_box=70,1178,496,1257>Age</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            144,
            145
        ],
        "focused": false,
        "bounds": [
            [
                70,
                1270
            ],
            [
                496,
                1380
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 141,
        "temp_id": 143,
        "size": "426*110",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "0687a7378dd71b5e288422535fee2f12",
        "bound_box": "70,1270,496,1380",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                70,
                1273
            ],
            [
                254,
                1333
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "26 years",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 143,
        "temp_id": 144,
        "size": "184*60",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]True[text]26 years[enabled,,]",
        "view_str": "4a6acc2906083a4816e2d968d9500efa",
        "bound_box": "70,1273,254,1333",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "54",
        "full_desc": "<button bound_box=70,1273,254,1333>26 years</button>",
        "desc": "<button bound_box=70,1273,254,1333>26 years</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                70,
                1330
            ],
            [
                496,
                1380
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "September 4, 1998",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 143,
        "temp_id": 145,
        "size": "426*50",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]September 4, 1998[enabled,,]",
        "view_str": "e98177e1a03b53cfc09ad6df0dccdd7d",
        "bound_box": "70,1330,496,1380",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "55",
        "full_desc": "<button bound_box=70,1330,496,1380>September 4, 1998</button>",
        "desc": "<button bound_box=70,1330,496,1380>September 4, 1998</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            147
        ],
        "focused": false,
        "bounds": [
            [
                553,
                1149
            ],
            [
                1042,
                1412
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 137,
        "temp_id": 146,
        "size": "489*263",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "ac94a2d925c06296926fff54f0722688",
        "bound_box": "553,1149,1042,1412",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            148
        ],
        "focused": false,
        "bounds": [
            [
                553,
                1149
            ],
            [
                1042,
                1412
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 146,
        "temp_id": 147,
        "size": "489*263",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "b3c93da92561da202820b96b91595908",
        "bound_box": "553,1149,1042,1412",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "56",
        "full_desc": "<button bound_box=553,1149,1042,1412></button>",
        "desc": "<button bound_box=553,1149,1042,1412></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            149,
            150
        ],
        "focused": false,
        "bounds": [
            [
                553,
                1149
            ],
            [
                1042,
                1412
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 147,
        "temp_id": 148,
        "size": "489*263",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "d716309c101c585822ca2c0b7bcb215f",
        "bound_box": "553,1149,1042,1412",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                588,
                1178
            ],
            [
                1010,
                1252
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_50",
        "checked": false,
        "text": "Founders",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 148,
        "temp_id": 149,
        "size": "422*74",
        "signature": "[class]android.widget.Button[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_50[visible]True[text]Founders[enabled,,]",
        "view_str": "71a48942da8f8bc371b77ce431c369e4",
        "bound_box": "588,1178,1010,1252",
        "content_free_signature": "[class]android.widget.Button[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_50[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "57",
        "full_desc": "<button bound_box=588,1178,1010,1252>Founders</button>",
        "desc": "<button bound_box=588,1178,1010,1252>Founders</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 3,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            151,
            153,
            155
        ],
        "focused": false,
        "bounds": [
            [
                588,
                1249
            ],
            [
                1010,
                1380
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 148,
        "temp_id": 150,
        "size": "422*131",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "42a4c8fbb953ac042e2d1a78efcce489",
        "bound_box": "588,1249,1010,1380",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            152
        ],
        "focused": false,
        "bounds": [
            [
                588,
                1288
            ],
            [
                874,
                1380
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 150,
        "temp_id": 151,
        "size": "286*92",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "b4f26bc0de21f381b6bbf78e5dd5bc0e",
        "bound_box": "588,1288,874,1380",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                588,
                1288
            ],
            [
                874,
                1380
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Larry Page, Sergey Brin",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 151,
        "temp_id": 152,
        "size": "286*92",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]Larry Page, Sergey Brin[enabled,,]",
        "view_str": "4382f893e3b7081f7b3177ef8ae58133",
        "bound_box": "588,1288,874,1380",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "58",
        "full_desc": "<button bound_box=588,1288,874,1380>Larry Page, Sergey Brin</button>",
        "desc": "<button bound_box=588,1288,874,1380>Larry Page, Sergey Brin</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            154
        ],
        "focused": false,
        "bounds": [
            [
                882,
                1249
            ],
            [
                1000,
                1367
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 150,
        "temp_id": 153,
        "size": "118*118",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "36774c20f1d15daac1d70f34fc084277",
        "bound_box": "882,1249,1000,1367",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                882,
                1249
            ],
            [
                1000,
                1367
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 153,
        "temp_id": 154,
        "size": "118*118",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "a5fc223c8bc05861263aaba3c68feaab",
        "bound_box": "882,1249,1000,1367",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            156
        ],
        "focused": false,
        "bounds": [
            [
                590,
                1333
            ],
            [
                1013,
                1396
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 150,
        "temp_id": 155,
        "size": "423*63",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "65a71fcfe6c3f65de2581ec6bb630232",
        "bound_box": "590,1333,1013,1396",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                939,
                1333
            ],
            [
                1013,
                1386
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "+1",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 155,
        "temp_id": 156,
        "size": "74*53",
        "signature": "[class]android.widget.Button[resource_id]None[visible]True[text]+1[enabled,,]",
        "view_str": "cc0f74a7119a3a34789e9ac06db28e29",
        "bound_box": "939,1333,1013,1386",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "59",
        "full_desc": "<button bound_box=939,1333,1013,1386>+1</button>",
        "desc": "<button bound_box=939,1333,1013,1386>+1</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                1451
            ],
            [
                1084,
                1522
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "See also",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 125,
        "temp_id": 157,
        "size": "1084*71",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]See also[enabled,,]",
        "view_str": "aa202903d36baff5cd54b0df3469645f",
        "bound_box": "0,1451,1084,1522",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "60",
        "full_desc": "<button bound_box=0,1451,1084,1522>See also</button>",
        "desc": "<button bound_box=0,1451,1084,1522>See also</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            159
        ],
        "focused": false,
        "bounds": [
            [
                0,
                1519
            ],
            [
                1084,
                1685
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 125,
        "temp_id": 158,
        "size": "1084*166",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "0360dc24dfa46471c7f1035e05465f8f",
        "bound_box": "0,1519,1084,1685",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            160
        ],
        "focused": false,
        "bounds": [
            [
                0,
                1519
            ],
            [
                1084,
                1685
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": true,
        "selected": false,
        "long_clickable": false,
        "parent": 158,
        "temp_id": 159,
        "size": "1084*166",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "a8d2be86fbd9b0241a81f1023bfe3ba2",
        "bound_box": "0,1519,1084,1685",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "scroll up",
            "scroll down",
            "scroll left",
            "scroll right"
        ],
        "status": [],
        "local_id": "61",
        "full_desc": "<button bound_box=0,1519,1084,1685></button>",
        "desc": "<button bound_box=0,1519,1084,1685></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 15,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            161,
            165,
            169,
            173,
            181,
            189,
            197,
            205,
            213
        ],
        "focused": false,
        "bounds": [
            [
                0,
                1519
            ],
            [
                5339,
                1685
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.widget.ListView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 159,
        "temp_id": 160,
        "size": "5339*166",
        "signature": "[class]android.widget.ListView[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "34a817f16255733cc562391f7f90292d",
        "bound_box": "0,1519,5339,1685",
        "content_free_signature": "[class]android.widget.ListView[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Apple",
        "children": [
            162,
            163
        ],
        "focused": false,
        "bounds": [
            [
                42,
                1519
            ],
            [
                343,
                1685
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 160,
        "temp_id": 161,
        "size": "301*166",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "097f1ee5336aa447a9d1d1905f0744eb",
        "bound_box": "42,1519,343,1685",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "62",
        "full_desc": "<button alt='Apple' bound_box=42,1519,343,1685></button>",
        "desc": "<button alt='Apple' bound_box=42,1519,343,1685></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                55,
                1538
            ],
            [
                186,
                1666
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 161,
        "temp_id": 162,
        "size": "131*128",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "146f75ae3778871bf47e0c6ea1c5acf7",
        "bound_box": "55,1538,186,1666",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            164
        ],
        "focused": false,
        "bounds": [
            [
                212,
                1577
            ],
            [
                312,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 161,
        "temp_id": 163,
        "size": "100*47",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "4ab6732377bc59dc20150d450e85fee5",
        "bound_box": "212,1577,312,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                212,
                1577
            ],
            [
                312,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Apple",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 163,
        "temp_id": 164,
        "size": "100*47",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]Apple[enabled,,]",
        "view_str": "921e5dc48d521b07c3c557789a45230b",
        "bound_box": "212,1577,312,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "63",
        "full_desc": "<button bound_box=212,1577,312,1624>Apple</button>",
        "desc": "<button bound_box=212,1577,312,1624>Apple</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Microsoft",
        "children": [
            166,
            167
        ],
        "focused": false,
        "bounds": [
            [
                370,
                1519
            ],
            [
                737,
                1685
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 160,
        "temp_id": 165,
        "size": "367*166",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "097f1ee5336aa447a9d1d1905f0744eb",
        "bound_box": "370,1519,737,1685",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "64",
        "full_desc": "<button alt='Microsoft' bound_box=370,1519,737,1685></button>",
        "desc": "<button alt='Microsoft' bound_box=370,1519,737,1685></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                385,
                1538
            ],
            [
                517,
                1666
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 165,
        "temp_id": 166,
        "size": "132*128",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "146f75ae3778871bf47e0c6ea1c5acf7",
        "bound_box": "385,1538,517,1666",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            168
        ],
        "focused": false,
        "bounds": [
            [
                543,
                1577
            ],
            [
                706,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 165,
        "temp_id": 167,
        "size": "163*47",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "44caf57868884d9b99ed3d0304be0a87",
        "bound_box": "543,1577,706,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                543,
                1577
            ],
            [
                706,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Microsoft",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 167,
        "temp_id": 168,
        "size": "163*47",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]Microsoft[enabled,,]",
        "view_str": "9b2cfa90f028160a212f71296574f968",
        "bound_box": "543,1577,706,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "65",
        "full_desc": "<button bound_box=543,1577,706,1624>Microsoft</button>",
        "desc": "<button bound_box=543,1577,706,1624>Microsoft</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Yelp",
        "children": [
            170,
            171
        ],
        "focused": false,
        "bounds": [
            [
                766,
                1519
            ],
            [
                1044,
                1685
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 160,
        "temp_id": 169,
        "size": "278*166",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "097f1ee5336aa447a9d1d1905f0744eb",
        "bound_box": "766,1519,1044,1685",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "66",
        "full_desc": "<button alt='Yelp' bound_box=766,1519,1044,1685></button>",
        "desc": "<button alt='Yelp' bound_box=766,1519,1044,1685></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                782,
                1538
            ],
            [
                910,
                1666
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 169,
        "temp_id": 170,
        "size": "128*128",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "146f75ae3778871bf47e0c6ea1c5acf7",
        "bound_box": "782,1538,910,1666",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            172
        ],
        "focused": false,
        "bounds": [
            [
                939,
                1577
            ],
            [
                1013,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 169,
        "temp_id": 171,
        "size": "74*47",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "f70078eaba01057268798772fcbe1b8e",
        "bound_box": "939,1577,1013,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                939,
                1577
            ],
            [
                1013,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Yelp",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 171,
        "temp_id": 172,
        "size": "74*47",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]Yelp[enabled,,]",
        "view_str": "746e75e785fa2746bce2614049b52e61",
        "bound_box": "939,1577,1013,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "67",
        "full_desc": "<button bound_box=939,1577,1013,1624>Yelp</button>",
        "desc": "<button bound_box=939,1577,1013,1624>Yelp</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Samsung Electronics",
        "children": [
            175
        ],
        "focused": false,
        "bounds": [
            [
                1073,
                1519
            ],
            [
                1614,
                1685
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_52",
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 160,
        "temp_id": 173,
        "size": "541*166",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_52[visible]True[text]None[enabled,,]",
        "view_str": "722b5eb1a253226525f7751986547529",
        "bound_box": "1073,1519,1614,1685",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_52[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "68",
        "full_desc": "<button alt='Samsung Electronics' bound_box=1073,1519,1614,1685></button>",
        "desc": "<button alt='Samsung Electronics' bound_box=1073,1519,1614,1685></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1089,
                1538
            ],
            [
                1218,
                1666
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 173,
        "temp_id": 174,
        "size": "129*128",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "b82fda2fd6c648e29b938f4859a2e890",
        "bound_box": "1089,1538,1218,1666",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            176
        ],
        "focused": false,
        "bounds": [
            [
                1246,
                1556
            ],
            [
                1582,
                1648
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 173,
        "temp_id": 175,
        "size": "336*92",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "e8479965e5791d111688304dcc1818cd",
        "bound_box": "1246,1556,1582,1648",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1246,
                1556
            ],
            [
                1582,
                1648
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Samsung Electronics",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 175,
        "temp_id": 176,
        "size": "336*92",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Samsung Electronics[enabled,,]",
        "view_str": "52eb6485a7f12ef71aaf99ca7b7d23c4",
        "bound_box": "1246,1556,1582,1648",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Altaba",
        "children": [
            178,
            179
        ],
        "focused": false,
        "bounds": [
            [
                1643,
                1519
            ],
            [
                1958,
                1685
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_56",
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 160,
        "temp_id": 177,
        "size": "315*166",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_56[visible]False[text]None[enabled,,]",
        "view_str": "84bc01e3b689a5bc59fd3d83d41421dd",
        "bound_box": "1643,1519,1958,1685",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_56[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1659,
                1538
            ],
            [
                1787,
                1666
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 177,
        "temp_id": 178,
        "size": "128*128",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "14057c549fd1e0d4596c0b9d116b5d58",
        "bound_box": "1659,1538,1787,1666",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            180
        ],
        "focused": false,
        "bounds": [
            [
                1816,
                1577
            ],
            [
                1926,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 177,
        "temp_id": 179,
        "size": "110*47",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "e9d106f7279a4b9a49f977b5d661e462",
        "bound_box": "1816,1577,1926,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1816,
                1577
            ],
            [
                1926,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Altaba",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 179,
        "temp_id": 180,
        "size": "110*47",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Altaba[enabled,,]",
        "view_str": "96cbb0c51a6617732146658edf40c471",
        "bound_box": "1816,1577,1926,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "YouTube",
        "children": [
            182,
            183
        ],
        "focused": false,
        "bounds": [
            [
                1984,
                1519
            ],
            [
                2338,
                1685
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_62",
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 160,
        "temp_id": 181,
        "size": "354*166",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_62[visible]False[text]None[enabled,,]",
        "view_str": "676aa7d29198a64ac0cf66006b771024",
        "bound_box": "1984,1519,2338,1685",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_62[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                2002,
                1538
            ],
            [
                2131,
                1666
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 181,
        "temp_id": 182,
        "size": "129*128",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "feac1172af5e9f687ac209e93fb7892d",
        "bound_box": "2002,1538,2131,1666",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            184
        ],
        "focused": false,
        "bounds": [
            [
                2157,
                1577
            ],
            [
                2307,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 181,
        "temp_id": 183,
        "size": "150*47",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "ab204f36132deecb19a890f3cbad2b21",
        "bound_box": "2157,1577,2307,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                2157,
                1577
            ],
            [
                2307,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "YouTube",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 183,
        "temp_id": 184,
        "size": "150*47",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]YouTube[enabled,,]",
        "view_str": "8f898d6d8e169052bc23e056aa7a1a82",
        "bound_box": "2157,1577,2307,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Meta",
        "children": [
            186,
            187
        ],
        "focused": false,
        "bounds": [
            [
                2365,
                1519
            ],
            [
                2659,
                1685
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_64",
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 160,
        "temp_id": 185,
        "size": "294*166",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_64[visible]False[text]None[enabled,,]",
        "view_str": "76512f39222fc732901e2ae05e513f57",
        "bound_box": "2365,1519,2659,1685",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_64[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                2380,
                1538
            ],
            [
                2512,
                1666
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 185,
        "temp_id": 186,
        "size": "132*128",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "2c3f8bac4ee7f5319dddd8084590c796",
        "bound_box": "2380,1538,2512,1666",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            188
        ],
        "focused": false,
        "bounds": [
            [
                2541,
                1577
            ],
            [
                2625,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 185,
        "temp_id": 187,
        "size": "84*47",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "8de48367144a2281a19cbf5f95276600",
        "bound_box": "2541,1577,2625,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                2541,
                1577
            ],
            [
                2625,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Meta",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 187,
        "temp_id": 188,
        "size": "84*47",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Meta[enabled,,]",
        "view_str": "23f4f2f342bf42e080a3986aa8aa48ea",
        "bound_box": "2541,1577,2625,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Canva",
        "children": [
            190,
            191
        ],
        "focused": false,
        "bounds": [
            [
                2685,
                1519
            ],
            [
                2995,
                1685
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_66",
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 160,
        "temp_id": 189,
        "size": "310*166",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_66[visible]False[text]None[enabled,,]",
        "view_str": "cdd86ab336025857d649a6c012759eba",
        "bound_box": "2685,1519,2995,1685",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_66[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                2701,
                1538
            ],
            [
                2832,
                1666
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 189,
        "temp_id": 190,
        "size": "131*128",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "af6a0d573f89074a512741799ee8994f",
        "bound_box": "2701,1538,2832,1666",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            192
        ],
        "focused": false,
        "bounds": [
            [
                2858,
                1577
            ],
            [
                2966,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 189,
        "temp_id": 191,
        "size": "108*47",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "9aa358f4644a8a7f228e856548408edc",
        "bound_box": "2858,1577,2966,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                2858,
                1577
            ],
            [
                2966,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Canva",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 191,
        "temp_id": 192,
        "size": "108*47",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Canva[enabled,,]",
        "view_str": "0ca19dc80d1a9468349c809aa5e77b18",
        "bound_box": "2858,1577,2966,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Baidu",
        "children": [
            194,
            195
        ],
        "focused": false,
        "bounds": [
            [
                3024,
                1519
            ],
            [
                3325,
                1685
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_68",
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 160,
        "temp_id": 193,
        "size": "301*166",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_68[visible]False[text]None[enabled,,]",
        "view_str": "35f572c9f09a6afc6782825e7d6c56bd",
        "bound_box": "3024,1519,3325,1685",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_68[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                3039,
                1538
            ],
            [
                3171,
                1666
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 193,
        "temp_id": 194,
        "size": "132*128",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "d6cf223f0d4d4cebd19874679fdaa639",
        "bound_box": "3039,1538,3171,1666",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            196
        ],
        "focused": false,
        "bounds": [
            [
                3197,
                1577
            ],
            [
                3294,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 193,
        "temp_id": 195,
        "size": "97*47",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "de451d332b65d958ca776fa1b0fb9d4f",
        "bound_box": "3197,1577,3294,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                3197,
                1577
            ],
            [
                3294,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Baidu",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 195,
        "temp_id": 196,
        "size": "97*47",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Baidu[enabled,,]",
        "view_str": "24f55b2fd0659d8f3b2ab2dd040cb937",
        "bound_box": "3197,1577,3294,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Amazon Web Services",
        "children": [
            198,
            199
        ],
        "focused": false,
        "bounds": [
            [
                3354,
                1519
            ],
            [
                3895,
                1685
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_70",
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 160,
        "temp_id": 197,
        "size": "541*166",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_70[visible]False[text]None[enabled,,]",
        "view_str": "ccbb4935ef82a53fb01d9d2087512d25",
        "bound_box": "3354,1519,3895,1685",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_70[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                3370,
                1538
            ],
            [
                3499,
                1666
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 197,
        "temp_id": 198,
        "size": "129*128",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "577759488e07651b19b3dea24589145d",
        "bound_box": "3370,1538,3499,1666",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            200
        ],
        "focused": false,
        "bounds": [
            [
                3528,
                1556
            ],
            [
                3864,
                1648
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 197,
        "temp_id": 199,
        "size": "336*92",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "ffc071f1cbbde6a8ba2c0a37e817902b",
        "bound_box": "3528,1556,3864,1648",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                3528,
                1556
            ],
            [
                3864,
                1648
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Amazon Web Services",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 199,
        "temp_id": 200,
        "size": "336*92",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Amazon Web Services[enabled,,]",
        "view_str": "4d199843eb478bb3ecab25fe26a911fd",
        "bound_box": "3528,1556,3864,1648",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "OpenAI",
        "children": [
            202,
            203
        ],
        "focused": false,
        "bounds": [
            [
                3924,
                1519
            ],
            [
                4252,
                1685
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_72",
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 160,
        "temp_id": 201,
        "size": "328*166",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_72[visible]False[text]None[enabled,,]",
        "view_str": "9be2478d658fbd27cb20d53a3a5467ed",
        "bound_box": "3924,1519,4252,1685",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_72[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                3940,
                1538
            ],
            [
                4068,
                1666
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 201,
        "temp_id": 202,
        "size": "128*128",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "19a4cc1283166b74edb85b6b517484e0",
        "bound_box": "3940,1538,4068,1666",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            204
        ],
        "focused": false,
        "bounds": [
            [
                4097,
                1577
            ],
            [
                4221,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 201,
        "temp_id": 203,
        "size": "124*47",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "c729638a0de0509db92f37dfbe55c897",
        "bound_box": "4097,1577,4221,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                4097,
                1577
            ],
            [
                4221,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "OpenAI",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 203,
        "temp_id": 204,
        "size": "124*47",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]OpenAI[enabled,,]",
        "view_str": "b3f3da16ac291101bb411c7282470a5a",
        "bound_box": "4097,1577,4221,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Netflix",
        "children": [
            206,
            207
        ],
        "focused": false,
        "bounds": [
            [
                4281,
                1519
            ],
            [
                4596,
                1685
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_74",
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 160,
        "temp_id": 205,
        "size": "315*166",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_74[visible]False[text]None[enabled,,]",
        "view_str": "bef67802f1ba8fbf90cf33b5f4c8022a",
        "bound_box": "4281,1519,4596,1685",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_74[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                4297,
                1538
            ],
            [
                4425,
                1666
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 205,
        "temp_id": 206,
        "size": "128*128",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "8b71e873eac2924bff3297b94dc98a53",
        "bound_box": "4297,1538,4425,1666",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            208
        ],
        "focused": false,
        "bounds": [
            [
                4454,
                1577
            ],
            [
                4564,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 205,
        "temp_id": 207,
        "size": "110*47",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "a8742e119380a2ed1b1709bec2967951",
        "bound_box": "4454,1577,4564,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                4454,
                1577
            ],
            [
                4564,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Netflix",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 207,
        "temp_id": 208,
        "size": "110*47",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Netflix[enabled,,]",
        "view_str": "f77ced66c6d135656b52d8adc5565f56",
        "bound_box": "4454,1577,4564,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Nvidia",
        "children": [
            210,
            211
        ],
        "focused": false,
        "bounds": [
            [
                4625,
                1519
            ],
            [
                4937,
                1685
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_76",
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 160,
        "temp_id": 209,
        "size": "312*166",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_76[visible]False[text]None[enabled,,]",
        "view_str": "64dafb29fdd91b389a7848daf101c1af",
        "bound_box": "4625,1519,4937,1685",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_76[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                4641,
                1538
            ],
            [
                4769,
                1666
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 209,
        "temp_id": 210,
        "size": "128*128",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "f4f8a65c495e8e6730e587c2e5d418f2",
        "bound_box": "4641,1538,4769,1666",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            212
        ],
        "focused": false,
        "bounds": [
            [
                4798,
                1577
            ],
            [
                4906,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 209,
        "temp_id": 211,
        "size": "108*47",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "3db3fbc0f09b290cc43b19545effb961",
        "bound_box": "4798,1577,4906,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                4798,
                1577
            ],
            [
                4906,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Nvidia",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 211,
        "temp_id": 212,
        "size": "108*47",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Nvidia[enabled,,]",
        "view_str": "e4be433f624ae0fb014103252a4cfd21",
        "bound_box": "4798,1577,4906,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Spotify",
        "children": [
            214,
            215
        ],
        "focused": false,
        "bounds": [
            [
                4963,
                1519
            ],
            [
                5289,
                1685
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_78",
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 160,
        "temp_id": 213,
        "size": "326*166",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_78[visible]False[text]None[enabled,,]",
        "view_str": "2393643f2084eae7cade08e1daf281e4",
        "bound_box": "4963,1519,5289,1685",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_78[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                4979,
                1538
            ],
            [
                5110,
                1666
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 213,
        "temp_id": 214,
        "size": "131*128",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "75d0372ab7f5bfb1517cee48173cfee9",
        "bound_box": "4979,1538,5110,1666",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            216
        ],
        "focused": false,
        "bounds": [
            [
                5137,
                1577
            ],
            [
                5257,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 213,
        "temp_id": 215,
        "size": "120*47",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "30caac877c092c3be908f5643db8f71d",
        "bound_box": "5137,1577,5257,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                5137,
                1577
            ],
            [
                5257,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Spotify",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 215,
        "temp_id": 216,
        "size": "120*47",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Spotify[enabled,,]",
        "view_str": "85f7ed94c7b43811c16be427b8de617a",
        "bound_box": "5137,1577,5257,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "GitHub",
        "children": [
            218,
            219
        ],
        "focused": false,
        "bounds": [
            [
                5318,
                1519
            ],
            [
                5638,
                1685
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_80",
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 160,
        "temp_id": 217,
        "size": "320*166",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_80[visible]False[text]None[enabled,,]",
        "view_str": "6cecc58552991f71fc02aee332d5f342",
        "bound_box": "5318,1519,5638,1685",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_80[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                5334,
                1538
            ],
            [
                5462,
                1666
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 217,
        "temp_id": 218,
        "size": "128*128",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "1027d8a3a2e0a2d6f60723ca8b399176",
        "bound_box": "5334,1538,5462,1666",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            220
        ],
        "focused": false,
        "bounds": [
            [
                5491,
                1577
            ],
            [
                5607,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 217,
        "temp_id": 219,
        "size": "116*47",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "58132b61a51b2bafe1eeca715a398bb2",
        "bound_box": "5491,1577,5607,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                5491,
                1577
            ],
            [
                5607,
                1624
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "GitHub",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 219,
        "temp_id": 220,
        "size": "116*47",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]GitHub[enabled,,]",
        "view_str": "4c145fa7b0f6b784fa8d64f7d5e791b4",
        "bound_box": "5491,1577,5607,1624",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                1748
            ],
            [
                1084,
                2026
            ]
        ],
        "resource_id": "fld_2-0yZ-jtAcyGptQPofi-iA8_2",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 123,
        "temp_id": 221,
        "size": "1084*278",
        "signature": "[class]android.view.View[resource_id]fld_2-0yZ-jtAcyGptQPofi-iA8_2[visible]True[text][enabled,,]",
        "view_str": "2c3c844c4372625871adf3562b3d54a6",
        "bound_box": "0,1748,1084,2026",
        "content_free_signature": "[class]android.view.View[resource_id]fld_2-0yZ-jtAcyGptQPofi-iA8_2[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            223,
            225
        ],
        "focused": false,
        "bounds": [
            [
                0,
                1748
            ],
            [
                1084,
                2026
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 123,
        "temp_id": 222,
        "size": "1084*278",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "a5ea6249ac66b430bc5b5aab55ccdfb1",
        "bound_box": "0,1748,1084,2026",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "69",
        "full_desc": "<button bound_box=0,1748,1084,2026></button>",
        "desc": "<button bound_box=0,1748,1084,2026></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            224
        ],
        "focused": false,
        "bounds": [
            [
                0,
                1748
            ],
            [
                225,
                1903
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 222,
        "temp_id": 223,
        "size": "225*155",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "799adb25945fb5b3177b35cbe117fe3b",
        "bound_box": "0,1748,225,1903",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                1790
            ],
            [
                183,
                1861
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "About",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 223,
        "temp_id": 224,
        "size": "141*71",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]About[enabled,,]",
        "view_str": "37f90ba78b9b0885d75b7f0545d3b465",
        "bound_box": "42,1790,183,1861",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "70",
        "full_desc": "<button bound_box=42,1790,183,1861>About</button>",
        "desc": "<button bound_box=42,1790,183,1861>About</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            226
        ],
        "focused": false,
        "bounds": [
            [
                0,
                1900
            ],
            [
                1084,
                1997
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 222,
        "temp_id": 225,
        "size": "1084*97",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "0360dc24dfa46471c7f1035e05465f8f",
        "bound_box": "0,1900,1084,1997",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "71",
        "full_desc": "<button bound_box=0,1900,1084,1997></button>",
        "desc": "<button bound_box=0,1900,1084,1997></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            227
        ],
        "focused": false,
        "bounds": [
            [
                42,
                1900
            ],
            [
                1042,
                1997
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 225,
        "temp_id": 226,
        "size": "1000*97",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "364a03bda94d02136cd0d0934997f947",
        "bound_box": "42,1900,1042,1997",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "72",
        "full_desc": "<button bound_box=42,1900,1042,1997></button>",
        "desc": "<button bound_box=42,1900,1042,1997></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "google.com",
        "children": [
            228
        ],
        "focused": false,
        "bounds": [
            [
                42,
                1900
            ],
            [
                1042,
                1997
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 226,
        "temp_id": 227,
        "size": "1000*97",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "ad15df6391356a69563642925cd03428",
        "bound_box": "42,1900,1042,1997",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "73",
        "full_desc": "<button alt='google.com' bound_box=42,1900,1042,1997></button>",
        "desc": "<button alt='google.com' bound_box=42,1900,1042,1997></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            229
        ],
        "focused": false,
        "bounds": [
            [
                42,
                1900
            ],
            [
                1042,
                1997
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 227,
        "temp_id": 228,
        "size": "1000*97",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "a0de06db5b079378a148abac0f8c7d57",
        "bound_box": "42,1900,1042,1997",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                1900
            ],
            [
                380,
                1997
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "google.com",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 228,
        "temp_id": 229,
        "size": "338*97",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]google.com[enabled,,]",
        "view_str": "d539f58178e9bcf2e6e697c9f4fc543c",
        "bound_box": "42,1900,380,1997",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "74",
        "full_desc": "<button bound_box=42,1900,380,1997>google.com</button>",
        "desc": "<button bound_box=42,1900,380,1997>google.com</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google",
        "children": [
            231
        ],
        "focused": false,
        "bounds": [
            [
                0,
                2021
            ],
            [
                1084,
                2218
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 119,
        "temp_id": 230,
        "size": "1084*197",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]None[enabled,,]",
        "view_str": "7137ae2b7bcc58aafec2375452e49cfa",
        "bound_box": "0,2021,1084,2218",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "75",
        "full_desc": "<button alt='Google' bound_box=0,2021,1084,2218></button>",
        "desc": "<button alt='Google' bound_box=0,2021,1084,2218></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            232
        ],
        "focused": false,
        "bounds": [
            [
                0,
                2063
            ],
            [
                1084,
                2212
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 230,
        "temp_id": 231,
        "size": "1084*149",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "ddb7e4653885df36d62e903779532df8",
        "bound_box": "0,2063,1084,2212",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            233,
            234
        ],
        "focused": false,
        "bounds": [
            [
                42,
                2063
            ],
            [
                1042,
                2170
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 231,
        "temp_id": 232,
        "size": "1000*107",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "e4bec1248e893bb69f0d624c97b0334f",
        "bound_box": "42,2063,1042,2170",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                443,
                2092
            ],
            [
                564,
                2139
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 232,
        "temp_id": 233,
        "size": "121*47",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]True[text]Google[enabled,,]",
        "view_str": "cccbbdd92d9494c4317fe16fc6b47841",
        "bound_box": "443,2092,564,2139",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "76",
        "full_desc": "<button bound_box=443,2092,564,2139>Google</button>",
        "desc": "<button bound_box=443,2092,564,2139>Google</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                2063
            ],
            [
                1042,
                2170
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 232,
        "temp_id": 234,
        "size": "1000*107",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "ad534f821d5c87937440894b95fb27bd",
        "bound_box": "42,2063,1042,2170",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                2236
            ],
            [
                1084,
                2236
            ]
        ],
        "resource_id": "z9PoV",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 103,
        "temp_id": 235,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]z9PoV[visible]False[text][enabled,,]",
        "view_str": "e0f6c22460f02993cdc4aee81d7faeb7",
        "bound_box": "0,2236,1084,2236",
        "content_free_signature": "[class]android.view.View[resource_id]z9PoV[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                2236
            ],
            [
                1084,
                2236
            ]
        ],
        "resource_id": "fld_2-0yZ-jtAcyGptQPofi-iA8_3",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 103,
        "temp_id": 236,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]fld_2-0yZ-jtAcyGptQPofi-iA8_3[visible]False[text][enabled,,]",
        "view_str": "93674ac134364a7456c4bbdb08d00072",
        "bound_box": "0,2236,1084,2236",
        "content_free_signature": "[class]android.view.View[resource_id]fld_2-0yZ-jtAcyGptQPofi-iA8_3[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 3,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            238,
            261
        ],
        "focused": false,
        "bounds": [
            [
                0,
                2236
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 103,
        "temp_id": 237,
        "size": "1084*40",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "4408b3f0813e25775e5f14b6297ce426",
        "bound_box": "0,2236,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "77",
        "full_desc": "<button bound_box=0,2236,1084,2276></button>",
        "desc": "<button bound_box=0,2236,1084,2276></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 5,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            239,
            247,
            255
        ],
        "focused": false,
        "bounds": [
            [
                0,
                2236
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 237,
        "temp_id": 238,
        "size": "1084*40",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "384e8893a5fe5801a92b125e620e65e9",
        "bound_box": "0,2236,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "78",
        "full_desc": "<button bound_box=0,2236,1084,2276></button>",
        "desc": "<button bound_box=0,2236,1084,2276></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            240
        ],
        "focused": false,
        "bounds": [
            [
                0,
                2236
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 238,
        "temp_id": 239,
        "size": "1084*40",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "c959eeba891fddbe7d55fa0603a61efc",
        "bound_box": "0,2236,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "79",
        "full_desc": "<button bound_box=0,2236,1084,2276></button>",
        "desc": "<button bound_box=0,2236,1084,2276></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            241
        ],
        "focused": false,
        "bounds": [
            [
                0,
                2236
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 239,
        "temp_id": 240,
        "size": "1084*40",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text][enabled,,]",
        "view_str": "7775f4a6ad0cdb827c0cfda452ea010b",
        "bound_box": "0,2236,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            242
        ],
        "focused": false,
        "bounds": [
            [
                0,
                2236
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Phone number … Google customer service",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 240,
        "temp_id": 241,
        "size": "1084*40",
        "signature": "[class]android.view.View[resource_id]None[visible]True[text]Phone number … Google customer service[enabled,,]",
        "view_str": "fa494e5a52d72fc7c7768a0847452870",
        "bound_box": "0,2236,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "80",
        "full_desc": "<button bound_box=0,2236,1084,2276>Phone number … Google customer service</button>",
        "desc": "<button bound_box=0,2236,1084,2276>Phone number … Google customer service</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                2236
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Phone number … Google customer service",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 241,
        "temp_id": 242,
        "size": "1084*40",
        "signature": "[class]android.widget.Button[resource_id]None[visible]True[text]Phone number … Google customer service[enabled,,]",
        "view_str": "dc8157a9f44cee19d617b92ab38c71aa",
        "bound_box": "0,2236,1084,2276",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "81",
        "full_desc": "<button bound_box=0,2236,1084,2276>Phone number … Google customer service</button>",
        "desc": "<button bound_box=0,2236,1084,2276>Phone number … Google customer service</button>"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            244
        ],
        "focused": false,
        "bounds": [
            [
                0,
                2443
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 238,
        "temp_id": 243,
        "size": "1084*-167",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "95c02557e7b301a03e89e20c067252fa",
        "bound_box": "0,2443,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            245
        ],
        "focused": false,
        "bounds": [
            [
                0,
                2443
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 243,
        "temp_id": 244,
        "size": "1084*-167",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "74a0f6a98a0f338b90e247f5c32078c5",
        "bound_box": "0,2443,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            246
        ],
        "focused": false,
        "bounds": [
            [
                0,
                2446
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Cost … How much does it cost to meet Google?",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 244,
        "temp_id": 245,
        "size": "1084*-170",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Cost … How much does it cost to meet Google?[enabled,,]",
        "view_str": "b7ef418ce740244a47bea4fe6a8139ad",
        "bound_box": "0,2446,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                2446
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Cost … How much does it cost to meet Google?",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 245,
        "temp_id": 246,
        "size": "1084*-170",
        "signature": "[class]android.widget.Button[resource_id]None[visible]False[text]Cost … How much does it cost to meet Google?[enabled,,]",
        "view_str": "715c7af54c91f3b9be476ee8501472a5",
        "bound_box": "0,2446,1084,2276",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            248
        ],
        "focused": false,
        "bounds": [
            [
                0,
                2656
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 238,
        "temp_id": 247,
        "size": "1084*-380",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "95c02557e7b301a03e89e20c067252fa",
        "bound_box": "0,2656,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            249
        ],
        "focused": false,
        "bounds": [
            [
                0,
                2656
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 247,
        "temp_id": 248,
        "size": "1084*-380",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "42ffcc397ae4f686e2cff4b80c064ded",
        "bound_box": "0,2656,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            250
        ],
        "focused": false,
        "bounds": [
            [
                0,
                2659
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Search … How to search with google",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 248,
        "temp_id": 249,
        "size": "1084*-383",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Search … How to search with google[enabled,,]",
        "view_str": "2b50fb5d8186eda5c50c0954b131f091",
        "bound_box": "0,2659,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                2659
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Search … How to search with google",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 249,
        "temp_id": 250,
        "size": "1084*-383",
        "signature": "[class]android.widget.Button[resource_id]None[visible]False[text]Search … How to search with google[enabled,,]",
        "view_str": "3f38151a26b42bdf03180684eeac0f44",
        "bound_box": "0,2659,1084,2276",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            252
        ],
        "focused": false,
        "bounds": [
            [
                0,
                2869
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 238,
        "temp_id": 251,
        "size": "1084*-593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "95c02557e7b301a03e89e20c067252fa",
        "bound_box": "0,2869,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            253
        ],
        "focused": false,
        "bounds": [
            [
                0,
                2869
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 251,
        "temp_id": 252,
        "size": "1084*-593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "7a079a6e6faeb60ebbb3224816891cf9",
        "bound_box": "0,2869,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            254
        ],
        "focused": false,
        "bounds": [
            [
                0,
                2871
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "History … Google history",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 252,
        "temp_id": 253,
        "size": "1084*-595",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]History … Google history[enabled,,]",
        "view_str": "1d6d772c3bf7e63431c36589ab245e35",
        "bound_box": "0,2871,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                2871
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "History … Google history",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 253,
        "temp_id": 254,
        "size": "1084*-595",
        "signature": "[class]android.widget.Button[resource_id]None[visible]False[text]History … Google history[enabled,,]",
        "view_str": "75a57754220e310616d5b167c165efb5",
        "bound_box": "0,2871,1084,2276",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            256
        ],
        "focused": false,
        "bounds": [
            [
                0,
                3081
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 238,
        "temp_id": 255,
        "size": "1084*-805",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "95c02557e7b301a03e89e20c067252fa",
        "bound_box": "0,3081,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            257
        ],
        "focused": false,
        "bounds": [
            [
                0,
                3081
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 255,
        "temp_id": 256,
        "size": "1084*-805",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "a99b04e5ee1993c03b12365375530156",
        "bound_box": "0,3081,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            258
        ],
        "focused": false,
        "bounds": [
            [
                0,
                3081
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Message … Message by google",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 256,
        "temp_id": 257,
        "size": "1084*-805",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Message … Message by google[enabled,,]",
        "view_str": "ebfcea3c25587d06ea872e47c74fa186",
        "bound_box": "0,3081,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                3081
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Message … Message by google",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 257,
        "temp_id": 258,
        "size": "1084*-805",
        "signature": "[class]android.widget.Button[resource_id]None[visible]False[text]Message … Message by google[enabled,,]",
        "view_str": "a524fdadb29cb71edafcc564b6883781",
        "bound_box": "0,3081,1084,2276",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            260
        ],
        "focused": false,
        "bounds": [
            [
                0,
                3577
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_106",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 237,
        "temp_id": 259,
        "size": "1084*-1301",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_106[visible]False[text][enabled,,]",
        "view_str": "00e09e5f38783b783e635680e0ba3ff9",
        "bound_box": "0,3577,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_106[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                3291
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_109",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 259,
        "temp_id": 260,
        "size": "1084*-1015",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_109[visible]False[text][enabled,,]",
        "view_str": "7c05e9bf8b30e71036441dbf5e71efa2",
        "bound_box": "0,3291,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_109[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                918,
                3304
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Feedback",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 237,
        "temp_id": 261,
        "size": "124*-1028",
        "signature": "[class]android.widget.Button[resource_id]None[visible]False[text]Feedback[enabled,,]",
        "view_str": "177de98f14f3ebdd564bc80e3889f465",
        "bound_box": "918,3304,1042,2276",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 3,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            263,
            264,
            275
        ],
        "focused": false,
        "bounds": [
            [
                0,
                3391
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 103,
        "temp_id": 262,
        "size": "1084*-1115",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "f0da66a844fc6e6637674b19436cf8ec",
        "bound_box": "0,3391,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                3391
            ],
            [
                5,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Web Result with Site Links",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 262,
        "temp_id": 263,
        "size": "5*-1115",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Web Result with Site Links[enabled,,]",
        "view_str": "609ab553db61b712506fc7a80d096dd3",
        "bound_box": "0,3391,5,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            265,
            273
        ],
        "focused": false,
        "bounds": [
            [
                0,
                3391
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 262,
        "temp_id": 264,
        "size": "1084*-1115",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "a539b7de1efdd6418174853bacbbcbb3",
        "bound_box": "0,3391,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            266,
            272
        ],
        "focused": false,
        "bounds": [
            [
                0,
                3391
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 264,
        "temp_id": 265,
        "size": "1084*-1115",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "e4b7a5645a408c07747884a42b1c3607",
        "bound_box": "0,3391,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google https://www.google.com Google",
        "children": [
            267,
            271
        ],
        "focused": false,
        "bounds": [
            [
                0,
                3391
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 265,
        "temp_id": 266,
        "size": "1084*-1115",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "f2ecec12496874c75e383504bc2b2194",
        "bound_box": "0,3391,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            268
        ],
        "focused": false,
        "bounds": [
            [
                42,
                3430
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 266,
        "temp_id": 267,
        "size": "1000*-1154",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "3ffb465ae073c922ed968e04e0c2c9fb",
        "bound_box": "42,3430,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            269,
            270
        ],
        "focused": false,
        "bounds": [
            [
                42,
                3430
            ],
            [
                937,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 267,
        "temp_id": 268,
        "size": "895*-1154",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "3007d12b206bb35c788b5ce0df8591e2",
        "bound_box": "42,3430,937,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                147,
                3433
            ],
            [
                501,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 268,
        "temp_id": 269,
        "size": "354*-1157",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Google[enabled,,]",
        "view_str": "69272f8849b83eb776737811c7a132bf",
        "bound_box": "147,3433,501,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                147,
                3488
            ],
            [
                501,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "https://www.google.com",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 268,
        "temp_id": 270,
        "size": "354*-1212",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]https://www.google.com[enabled,,]",
        "view_str": "34c742875316ccedeabe30c9cba3931b",
        "bound_box": "147,3488,501,2276",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                3559
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 266,
        "temp_id": 271,
        "size": "1000*-1283",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Google[enabled,,]",
        "view_str": "4cef01b6966b79216e9d4eec027ad2c1",
        "bound_box": "42,3559,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                952,
                3391
            ],
            [
                1081,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "About this result",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 265,
        "temp_id": 272,
        "size": "129*-1115",
        "signature": "[class]android.widget.Button[resource_id]None[visible]False[text]About this result[enabled,,]",
        "view_str": "f001a46fdc92fe2611f7d32e0bdf4ef8",
        "bound_box": "952,3391,1081,2276",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            274
        ],
        "focused": false,
        "bounds": [
            [
                0,
                3617
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "tsuid_2-0yZ-jtAcyGptQPofi-iA8_128",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 264,
        "temp_id": 273,
        "size": "1084*-1341",
        "signature": "[class]android.view.View[resource_id]tsuid_2-0yZ-jtAcyGptQPofi-iA8_128[visible]False[text][enabled,,]",
        "view_str": "75a790ad048838eda92b0667b5080c0b",
        "bound_box": "0,3617,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]tsuid_2-0yZ-jtAcyGptQPofi-iA8_128[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                3648
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Search the world's information, including webpages, images, videos and more. Google has many special features to help you find exactly what you're looking ...",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 273,
        "temp_id": 274,
        "size": "1000*-1372",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "997f54715041054db797ef4ae543db19",
        "bound_box": "42,3648,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 12,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            276,
            277,
            279,
            280,
            282,
            283,
            285,
            286,
            288,
            289,
            291,
            292
        ],
        "focused": false,
        "bounds": [
            [
                0,
                3835
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 262,
        "temp_id": 275,
        "size": "1084*-1559",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "1699769a6efeba7768d53213867ad50c",
        "bound_box": "0,3835,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                3835
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 275,
        "temp_id": 276,
        "size": "1000*-1559",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "347aa7e60c4112dc4f0f88951ac6c267",
        "bound_box": "42,3835,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Accounts",
        "children": [
            278
        ],
        "focused": false,
        "bounds": [
            [
                42,
                3837
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 275,
        "temp_id": 277,
        "size": "1000*-1561",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "1a954497a16c194d61c3562f61c99a7c",
        "bound_box": "42,3837,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                3879
            ],
            [
                947,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Accounts",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 277,
        "temp_id": 278,
        "size": "905*-1603",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Accounts[enabled,,]",
        "view_str": "be452d44f6a2e6ae89f71f86d8dfcda2",
        "bound_box": "42,3879,947,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                3990
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 275,
        "temp_id": 279,
        "size": "1000*-1714",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "347aa7e60c4112dc4f0f88951ac6c267",
        "bound_box": "42,3990,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Flights",
        "children": [
            281
        ],
        "focused": false,
        "bounds": [
            [
                42,
                3992
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 275,
        "temp_id": 280,
        "size": "1000*-1716",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "8beb3feee2b654fe3c77239a617995c1",
        "bound_box": "42,3992,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                4034
            ],
            [
                947,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Flights",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 280,
        "temp_id": 281,
        "size": "905*-1758",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Flights[enabled,,]",
        "view_str": "0921f3038cf5f0ff20cb7ac8ea5bc39f",
        "bound_box": "42,4034,947,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                4144
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 275,
        "temp_id": 282,
        "size": "1000*-1868",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "347aa7e60c4112dc4f0f88951ac6c267",
        "bound_box": "42,4144,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Sign in",
        "children": [
            284
        ],
        "focused": false,
        "bounds": [
            [
                42,
                4147
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 275,
        "temp_id": 283,
        "size": "1000*-1871",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "ea90da9ca7a9d9cfd5388e78256f37e0",
        "bound_box": "42,4147,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                4189
            ],
            [
                947,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Sign in",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 283,
        "temp_id": 284,
        "size": "905*-1913",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Sign in[enabled,,]",
        "view_str": "9bbe60e34ccb4c00bba0696eb0f2cf66",
        "bound_box": "42,4189,947,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                4299
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 275,
        "temp_id": 285,
        "size": "1000*-2023",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "347aa7e60c4112dc4f0f88951ac6c267",
        "bound_box": "42,4299,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Docs",
        "children": [
            287
        ],
        "focused": false,
        "bounds": [
            [
                42,
                4302
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 275,
        "temp_id": 286,
        "size": "1000*-2026",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "ffec205db7382f1b58ea1c92da542b5c",
        "bound_box": "42,4302,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                4344
            ],
            [
                947,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Docs",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 286,
        "temp_id": 287,
        "size": "905*-2068",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Docs[enabled,,]",
        "view_str": "757168de239af524c6e0522ac6f283f5",
        "bound_box": "42,4344,947,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                4454
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 275,
        "temp_id": 288,
        "size": "1000*-2178",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "347aa7e60c4112dc4f0f88951ac6c267",
        "bound_box": "42,4454,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Translate",
        "children": [
            290
        ],
        "focused": false,
        "bounds": [
            [
                42,
                4457
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 275,
        "temp_id": 289,
        "size": "1000*-2181",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "39efda7df5cd46b781591d7d841100e9",
        "bound_box": "42,4457,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                4499
            ],
            [
                947,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Translate",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 289,
        "temp_id": 290,
        "size": "905*-2223",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Translate[enabled,,]",
        "view_str": "76a214f1709c56882e1d5fed2cfe6273",
        "bound_box": "42,4499,947,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                4609
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 275,
        "temp_id": 291,
        "size": "1000*-2333",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "347aa7e60c4112dc4f0f88951ac6c267",
        "bound_box": "42,4609,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Scholar",
        "children": [
            293
        ],
        "focused": false,
        "bounds": [
            [
                42,
                4609
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 275,
        "temp_id": 292,
        "size": "1000*-2333",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "75feab7cae276c4496f1127f8d344cbd",
        "bound_box": "42,4609,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                4651
            ],
            [
                947,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Scholar",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 292,
        "temp_id": 293,
        "size": "905*-2375",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Scholar[enabled,,]",
        "view_str": "bb1f4d57b8b92aa7893ff41a78dbe766",
        "bound_box": "42,4651,947,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            295
        ],
        "focused": false,
        "bounds": [
            [
                0,
                4782
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 103,
        "temp_id": 294,
        "size": "1084*-2506",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "67049e768ef110aa9225cda8bf46cb44",
        "bound_box": "0,4782,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 4,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            296,
            297,
            298,
            299
        ],
        "focused": false,
        "bounds": [
            [
                0,
                4782
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 294,
        "temp_id": 295,
        "size": "1084*-2506",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "2ac4d2c8494f123b3c204178f6b2ef06",
        "bound_box": "0,4782,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                4782
            ],
            [
                1168,
                2276
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_89",
        "checked": false,
        "text": "Install Google Google Play Google Rated 4.5 out of 5, (27M)",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 295,
        "temp_id": 296,
        "size": "1168*-2506",
        "signature": "[class]android.widget.Button[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_89[visible]False[text]None[enabled,,]",
        "view_str": "2e41077388caf709342dcc9970eae0d4",
        "bound_box": "0,4782,1168,2276",
        "content_free_signature": "[class]android.widget.Button[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_89[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                952,
                4782
            ],
            [
                1081,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "About this result",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 295,
        "temp_id": 297,
        "size": "129*-2506",
        "signature": "[class]android.widget.Button[resource_id]None[visible]False[text]About this result[enabled,,]",
        "view_str": "ed81035357963f4343806ff5f22b6f50",
        "bound_box": "952,4782,1081,2276",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                5105
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_90",
        "checked": false,
        "text": "About this app. arrow_forward. The Google app keeps you in the know about things that matter to you. Find quick answers, explore your interests, and stay up to ...",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 295,
        "temp_id": 298,
        "size": "1000*-2829",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_90[visible]False[text]None[enabled,,]",
        "view_str": "e3131c0f2318b4a95bc14a8eabcbccd7",
        "bound_box": "42,5105,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_90[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            300
        ],
        "focused": false,
        "bounds": [
            [
                0,
                5281
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_91",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 295,
        "temp_id": 299,
        "size": "1084*-3005",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_91[visible]False[text][enabled,,]",
        "view_str": "cf1740989c9718d3907bc708ed9e955d",
        "bound_box": "0,5281,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_91[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            301
        ],
        "focused": false,
        "bounds": [
            [
                795,
                5281
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 299,
        "temp_id": 300,
        "size": "247*-3005",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "3d440eff8814d99fbf09b2fa3e864ab5",
        "bound_box": "795,5281,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                795,
                5281
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_93",
        "checked": false,
        "text": "Install Google",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 300,
        "temp_id": 301,
        "size": "247*-3005",
        "signature": "[class]android.widget.Button[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_93[visible]False[text]Install Google[enabled,,]",
        "view_str": "d4e7efe74d3a28642c26a0d79ff38023",
        "bound_box": "795,5281,1042,2276",
        "content_free_signature": "[class]android.widget.Button[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_93[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 17,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            303,
            304,
            305,
            306,
            309,
            362,
            363,
            368,
            369,
            374,
            375,
            380,
            381,
            386,
            387,
            392,
            393
        ],
        "focused": false,
        "bounds": [
            [
                0,
                5439
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 103,
        "temp_id": 302,
        "size": "1084*-3163",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "3c7ace5c1efaaa88806691a735020369",
        "bound_box": "0,5439,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                5439
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 302,
        "temp_id": 303,
        "size": "1084*-3163",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "1b8d777b897133b175242f53ed4a7a08",
        "bound_box": "0,5439,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                7016
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 302,
        "temp_id": 304,
        "size": "1084*-4740",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "1b8d777b897133b175242f53ed4a7a08",
        "bound_box": "0,7016,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                5439
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 302,
        "temp_id": 305,
        "size": "1084*-3163",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "1b8d777b897133b175242f53ed4a7a08",
        "bound_box": "0,5439,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            307,
            308
        ],
        "focused": false,
        "bounds": [
            [
                0,
                5439
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 302,
        "temp_id": 306,
        "size": "1084*-3163",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "0a48bc6bdccf4585335f4aebb8f76bce",
        "bound_box": "0,5439,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                5481
            ],
            [
                1010,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "People also search for",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 306,
        "temp_id": 307,
        "size": "968*-3205",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]People also search for[enabled,,]",
        "view_str": "0f290b340c7c6e21bd663202f21621d9",
        "bound_box": "42,5481,1010,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                952,
                5439
            ],
            [
                1081,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "About this result",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 306,
        "temp_id": 308,
        "size": "129*-3163",
        "signature": "[class]android.widget.Button[resource_id]None[visible]False[text]About this result[enabled,,]",
        "view_str": "ed81035357963f4343806ff5f22b6f50",
        "bound_box": "952,5439,1081,2276",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            310
        ],
        "focused": false,
        "bounds": [
            [
                0,
                5622
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_135",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 302,
        "temp_id": 309,
        "size": "1084*-3346",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_135[visible]False[text][enabled,,]",
        "view_str": "2fc57ca4fff96433debda690280f4b56",
        "bound_box": "0,5622,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_135[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            311
        ],
        "focused": false,
        "bounds": [
            [
                0,
                5622
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "2-0yZ-jtAcyGptQPofi-iA8__78",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 309,
        "temp_id": 310,
        "size": "1084*-3346",
        "signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__78[visible]False[text][enabled,,]",
        "view_str": "95c75eb9cdc109d2b7221ffff47287c3",
        "bound_box": "0,5622,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__78[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            312
        ],
        "focused": false,
        "bounds": [
            [
                0,
                5622
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 310,
        "temp_id": 311,
        "size": "1084*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "0192476dd01e636d30b8e07ab91903c6",
        "bound_box": "0,5622,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            313
        ],
        "focused": false,
        "bounds": [
            [
                0,
                5622
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 311,
        "temp_id": 312,
        "size": "1084*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "db545ee17e26245c1cb520bc696cd216",
        "bound_box": "0,5622,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            314
        ],
        "focused": false,
        "bounds": [
            [
                0,
                5622
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 312,
        "temp_id": 313,
        "size": "1084*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "07a2631a3cebc98868694f265d498445",
        "bound_box": "0,5622,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            315,
            361
        ],
        "focused": false,
        "bounds": [
            [
                0,
                5622
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 313,
        "temp_id": 314,
        "size": "1084*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "74651e19ff7cf168b861c5e48ca1b7c0",
        "bound_box": "0,5622,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            316
        ],
        "focused": false,
        "bounds": [
            [
                0,
                5622
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": true,
        "selected": false,
        "long_clickable": false,
        "parent": 314,
        "temp_id": 315,
        "size": "1084*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "db4fe59f6da08d85530d7c2668d52597",
        "bound_box": "0,5622,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 8,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            317,
            322,
            327,
            332,
            337,
            343,
            349,
            355
        ],
        "focused": false,
        "bounds": [
            [
                0,
                5622
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.widget.ListView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 315,
        "temp_id": 316,
        "size": "1084*-3346",
        "signature": "[class]android.widget.ListView[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "9d03b7a9f0c6992bf174d22ffc1c3a2e",
        "bound_box": "0,5622,1084,2276",
        "content_free_signature": "[class]android.widget.ListView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            318
        ],
        "focused": false,
        "bounds": [
            [
                0,
                5622
            ],
            [
                357,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 316,
        "temp_id": 317,
        "size": "357*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "2b840f7b28ccf38e818c41361b580c8a",
        "bound_box": "0,5622,357,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            319,
            320
        ],
        "focused": false,
        "bounds": [
            [
                42,
                5622
            ],
            [
                325,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 317,
        "temp_id": 318,
        "size": "283*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "77b83576e0684251d3134bdbd21488f6",
        "bound_box": "42,5622,325,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google Maps",
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                5622
            ],
            [
                325,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 318,
        "temp_id": 319,
        "size": "283*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "fd517d5f712c840ab0c751a871cbc32d",
        "bound_box": "42,5622,325,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            321
        ],
        "focused": false,
        "bounds": [
            [
                42,
                5622
            ],
            [
                325,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 318,
        "temp_id": 320,
        "size": "283*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "67cc427e87b57211081c8c7ef3b44efd",
        "bound_box": "42,5622,325,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                5622
            ],
            [
                325,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 320,
        "temp_id": 321,
        "size": "283*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "7a4322a42254f89261c1a7a1cb664a02",
        "bound_box": "42,5622,325,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            323
        ],
        "focused": false,
        "bounds": [
            [
                351,
                5622
            ],
            [
                669,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 316,
        "temp_id": 322,
        "size": "318*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "2b840f7b28ccf38e818c41361b580c8a",
        "bound_box": "351,5622,669,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            324,
            325
        ],
        "focused": false,
        "bounds": [
            [
                351,
                5622
            ],
            [
                637,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 322,
        "temp_id": 323,
        "size": "286*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "77b83576e0684251d3134bdbd21488f6",
        "bound_box": "351,5622,637,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google Search",
        "children": [],
        "focused": false,
        "bounds": [
            [
                351,
                5622
            ],
            [
                637,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 323,
        "temp_id": 324,
        "size": "286*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "fd517d5f712c840ab0c751a871cbc32d",
        "bound_box": "351,5622,637,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            326
        ],
        "focused": false,
        "bounds": [
            [
                351,
                5622
            ],
            [
                637,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 323,
        "temp_id": 325,
        "size": "286*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "67cc427e87b57211081c8c7ef3b44efd",
        "bound_box": "351,5622,637,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                351,
                5622
            ],
            [
                637,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 325,
        "temp_id": 326,
        "size": "286*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "7a4322a42254f89261c1a7a1cb664a02",
        "bound_box": "351,5622,637,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            328
        ],
        "focused": false,
        "bounds": [
            [
                666,
                5622
            ],
            [
                981,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 316,
        "temp_id": 327,
        "size": "315*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "2b840f7b28ccf38e818c41361b580c8a",
        "bound_box": "666,5622,981,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            329,
            330
        ],
        "focused": false,
        "bounds": [
            [
                666,
                5622
            ],
            [
                950,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 327,
        "temp_id": 328,
        "size": "284*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "77b83576e0684251d3134bdbd21488f6",
        "bound_box": "666,5622,950,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google Classroom",
        "children": [],
        "focused": false,
        "bounds": [
            [
                666,
                5622
            ],
            [
                950,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 328,
        "temp_id": 329,
        "size": "284*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "fd517d5f712c840ab0c751a871cbc32d",
        "bound_box": "666,5622,950,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            331
        ],
        "focused": false,
        "bounds": [
            [
                666,
                5622
            ],
            [
                950,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 328,
        "temp_id": 330,
        "size": "284*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "67cc427e87b57211081c8c7ef3b44efd",
        "bound_box": "666,5622,950,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                666,
                5622
            ],
            [
                950,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 330,
        "temp_id": 331,
        "size": "284*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "7a4322a42254f89261c1a7a1cb664a02",
        "bound_box": "666,5622,950,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            333
        ],
        "focused": false,
        "bounds": [
            [
                979,
                5622
            ],
            [
                1294,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 316,
        "temp_id": 332,
        "size": "315*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "2b840f7b28ccf38e818c41361b580c8a",
        "bound_box": "979,5622,1294,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            334,
            335
        ],
        "focused": false,
        "bounds": [
            [
                979,
                5622
            ],
            [
                1262,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 332,
        "temp_id": 333,
        "size": "283*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "77b83576e0684251d3134bdbd21488f6",
        "bound_box": "979,5622,1262,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Gmail",
        "children": [],
        "focused": false,
        "bounds": [
            [
                979,
                5622
            ],
            [
                1262,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 333,
        "temp_id": 334,
        "size": "283*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "fd517d5f712c840ab0c751a871cbc32d",
        "bound_box": "979,5622,1262,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            336
        ],
        "focused": false,
        "bounds": [
            [
                979,
                5622
            ],
            [
                1262,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 333,
        "temp_id": 335,
        "size": "283*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "67cc427e87b57211081c8c7ef3b44efd",
        "bound_box": "979,5622,1262,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                979,
                5622
            ],
            [
                1262,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 335,
        "temp_id": 336,
        "size": "283*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "7a4322a42254f89261c1a7a1cb664a02",
        "bound_box": "979,5622,1262,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            338
        ],
        "focused": false,
        "bounds": [
            [
                1291,
                5622
            ],
            [
                1609,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 316,
        "temp_id": 337,
        "size": "318*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "c0175cbe6336279f1b24eb7b915b76ca",
        "bound_box": "1291,5622,1609,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            339
        ],
        "focused": false,
        "bounds": [
            [
                1291,
                5622
            ],
            [
                1575,
                2276
            ]
        ],
        "resource_id": "tsuid_2-0yZ-jtAcyGptQPofi-iA8_125",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 337,
        "temp_id": 338,
        "size": "284*-3346",
        "signature": "[class]android.view.View[resource_id]tsuid_2-0yZ-jtAcyGptQPofi-iA8_125[visible]False[text][enabled,,]",
        "view_str": "191260de07a85db72c76d8bc7edeea61",
        "bound_box": "1291,5622,1575,2276",
        "content_free_signature": "[class]android.view.View[resource_id]tsuid_2-0yZ-jtAcyGptQPofi-iA8_125[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            340,
            341
        ],
        "focused": false,
        "bounds": [
            [
                1291,
                5622
            ],
            [
                1575,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 338,
        "temp_id": 339,
        "size": "284*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "3470cdbcf491e093db41d53e5354346a",
        "bound_box": "1291,5622,1575,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google Chrome",
        "children": [],
        "focused": false,
        "bounds": [
            [
                1291,
                5622
            ],
            [
                1575,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 339,
        "temp_id": 340,
        "size": "284*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "e6e050048eb06abcdad02a2eba521a0f",
        "bound_box": "1291,5622,1575,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            342
        ],
        "focused": false,
        "bounds": [
            [
                1291,
                5622
            ],
            [
                1575,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 339,
        "temp_id": 341,
        "size": "284*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "727900e52d5d5271ce2c241d46535409",
        "bound_box": "1291,5622,1575,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1291,
                5622
            ],
            [
                1575,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 341,
        "temp_id": 342,
        "size": "284*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "ed8c0d9d2b7c8c087d79168d7b3f5c52",
        "bound_box": "1291,5622,1575,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            344
        ],
        "focused": false,
        "bounds": [
            [
                1603,
                5622
            ],
            [
                1921,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 316,
        "temp_id": 343,
        "size": "318*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "8284fd48b19da755f581e2b7e7904ba5",
        "bound_box": "1603,5622,1921,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            345
        ],
        "focused": false,
        "bounds": [
            [
                1603,
                5622
            ],
            [
                1890,
                2276
            ]
        ],
        "resource_id": "tsuid_2-0yZ-jtAcyGptQPofi-iA8_129",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 343,
        "temp_id": 344,
        "size": "287*-3346",
        "signature": "[class]android.view.View[resource_id]tsuid_2-0yZ-jtAcyGptQPofi-iA8_129[visible]False[text][enabled,,]",
        "view_str": "6842b341b9a0b69f1ad0c27d8a3fee5c",
        "bound_box": "1603,5622,1890,2276",
        "content_free_signature": "[class]android.view.View[resource_id]tsuid_2-0yZ-jtAcyGptQPofi-iA8_129[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            346,
            347
        ],
        "focused": false,
        "bounds": [
            [
                1603,
                5622
            ],
            [
                1890,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 344,
        "temp_id": 345,
        "size": "287*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "bc0357740fb5b8c0548448d9c3f74ff9",
        "bound_box": "1603,5622,1890,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google",
        "children": [],
        "focused": false,
        "bounds": [
            [
                1603,
                5622
            ],
            [
                1890,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 345,
        "temp_id": 346,
        "size": "287*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "af1093b9fba86a6a2a75ca6062ad0498",
        "bound_box": "1603,5622,1890,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            348
        ],
        "focused": false,
        "bounds": [
            [
                1603,
                5622
            ],
            [
                1890,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 345,
        "temp_id": 347,
        "size": "287*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "f776f04b11f775c7c15d4b6bdf293550",
        "bound_box": "1603,5622,1890,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1603,
                5622
            ],
            [
                1890,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 347,
        "temp_id": 348,
        "size": "287*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "284b9231b06e5f15085246b600d0b16e",
        "bound_box": "1603,5622,1890,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            350
        ],
        "focused": false,
        "bounds": [
            [
                1916,
                5622
            ],
            [
                2233,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 316,
        "temp_id": 349,
        "size": "317*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "ce6c46df8ec481ec5fce96aa3548a9d4",
        "bound_box": "1916,5622,2233,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            351
        ],
        "focused": false,
        "bounds": [
            [
                1916,
                5622
            ],
            [
                2202,
                2276
            ]
        ],
        "resource_id": "tsuid_2-0yZ-jtAcyGptQPofi-iA8_132",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 349,
        "temp_id": 350,
        "size": "286*-3346",
        "signature": "[class]android.view.View[resource_id]tsuid_2-0yZ-jtAcyGptQPofi-iA8_132[visible]False[text][enabled,,]",
        "view_str": "fe06324ca442e4d8da378660ce427c41",
        "bound_box": "1916,5622,2202,2276",
        "content_free_signature": "[class]android.view.View[resource_id]tsuid_2-0yZ-jtAcyGptQPofi-iA8_132[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            352,
            353
        ],
        "focused": false,
        "bounds": [
            [
                1916,
                5622
            ],
            [
                2202,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 350,
        "temp_id": 351,
        "size": "286*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "d30b324ef52842e5fcbcb823167c3c86",
        "bound_box": "1916,5622,2202,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google Lens",
        "children": [],
        "focused": false,
        "bounds": [
            [
                1916,
                5622
            ],
            [
                2202,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 351,
        "temp_id": 352,
        "size": "286*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "e94bb98377122970ee590b03f8843b5b",
        "bound_box": "1916,5622,2202,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            354
        ],
        "focused": false,
        "bounds": [
            [
                1916,
                5622
            ],
            [
                2202,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 351,
        "temp_id": 353,
        "size": "286*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "e791b1ca7ec9c095af8e09ea7a0a80de",
        "bound_box": "1916,5622,2202,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1916,
                5622
            ],
            [
                2202,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 353,
        "temp_id": 354,
        "size": "286*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "ac7f6ab70fa1ccb79267c84954ec5411",
        "bound_box": "1916,5622,2202,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            356
        ],
        "focused": false,
        "bounds": [
            [
                2228,
                5622
            ],
            [
                2556,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 316,
        "temp_id": 355,
        "size": "328*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "7d09174dc47b8eeacae6f7e29a65a5af",
        "bound_box": "2228,5622,2556,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            357
        ],
        "focused": false,
        "bounds": [
            [
                2228,
                5622
            ],
            [
                2514,
                2276
            ]
        ],
        "resource_id": "tsuid_2-0yZ-jtAcyGptQPofi-iA8_142",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 355,
        "temp_id": 356,
        "size": "286*-3346",
        "signature": "[class]android.view.View[resource_id]tsuid_2-0yZ-jtAcyGptQPofi-iA8_142[visible]False[text][enabled,,]",
        "view_str": "ceee092eb03683ac4fd5ee465966e9ca",
        "bound_box": "2228,5622,2514,2276",
        "content_free_signature": "[class]android.view.View[resource_id]tsuid_2-0yZ-jtAcyGptQPofi-iA8_142[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            358,
            359
        ],
        "focused": false,
        "bounds": [
            [
                2228,
                5622
            ],
            [
                2514,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 356,
        "temp_id": 357,
        "size": "286*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "3d12c60a463d5abb7389bc01a593ad07",
        "bound_box": "2228,5622,2514,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google Sites",
        "children": [],
        "focused": false,
        "bounds": [
            [
                2228,
                5622
            ],
            [
                2514,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 357,
        "temp_id": 358,
        "size": "286*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "6a7ac70bc9a7b0ec746261030e3fa4f1",
        "bound_box": "2228,5622,2514,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            360
        ],
        "focused": false,
        "bounds": [
            [
                2228,
                5622
            ],
            [
                2514,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 357,
        "temp_id": 359,
        "size": "286*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "80f05d9d99544aa79380801a5503f5ee",
        "bound_box": "2228,5622,2514,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                2228,
                5622
            ],
            [
                2514,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 359,
        "temp_id": 360,
        "size": "286*-3346",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "1d70473bdfd1c0ae9a7c4f6ca03106f3",
        "bound_box": "2228,5622,2514,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                459,
                6050
            ],
            [
                622,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 314,
        "temp_id": 361,
        "size": "163*-3774",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "bfccf2b99d698bd81a27960b1726d202",
        "bound_box": "459,6050,622,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                6129
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 302,
        "temp_id": 362,
        "size": "1000*-3853",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "1b8d777b897133b175242f53ed4a7a08",
        "bound_box": "42,6129,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            364
        ],
        "focused": false,
        "bounds": [
            [
                42,
                6132
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": "2-0yZ-jtAcyGptQPofi-iA8__80",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 302,
        "temp_id": 363,
        "size": "1000*-3856",
        "signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__80[visible]False[text][enabled,,]",
        "view_str": "1f2c74052b5b981d88acbf570c4b8f4c",
        "bound_box": "42,6132,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__80[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            365
        ],
        "focused": false,
        "bounds": [
            [
                42,
                6132
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 363,
        "temp_id": 364,
        "size": "1000*-3856",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "9be48132e99c895b7317d9e63bba8341",
        "bound_box": "42,6132,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "www.google search web",
        "children": [
            366,
            367
        ],
        "focused": false,
        "bounds": [
            [
                42,
                6132
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 364,
        "temp_id": 365,
        "size": "1000*-3856",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "93b9c4f7c3c4a81fd90b73621272df22",
        "bound_box": "42,6132,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                6184
            ],
            [
                916,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "www.google search web",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 365,
        "temp_id": 366,
        "size": "874*-3908",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]www.google search web[enabled,,]",
        "view_str": "67963458c29331a54046bcffb2f9017d",
        "bound_box": "42,6184,916,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                968,
                6184
            ],
            [
                1023,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.widget.Image",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 365,
        "temp_id": 367,
        "size": "55*-3908",
        "signature": "[class]android.widget.Image[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "bfa411f43067a7d44131c3f73d312fad",
        "bound_box": "968,6184,1023,2276",
        "content_free_signature": "[class]android.widget.Image[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                6289
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 302,
        "temp_id": 368,
        "size": "1000*-4013",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "1b8d777b897133b175242f53ed4a7a08",
        "bound_box": "42,6289,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            370
        ],
        "focused": false,
        "bounds": [
            [
                42,
                6292
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": "2-0yZ-jtAcyGptQPofi-iA8__83",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 302,
        "temp_id": 369,
        "size": "1000*-4016",
        "signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__83[visible]False[text][enabled,,]",
        "view_str": "0852291c011d5a2aa09120aa3edd7237",
        "bound_box": "42,6292,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__83[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            371
        ],
        "focused": false,
        "bounds": [
            [
                42,
                6292
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 369,
        "temp_id": 370,
        "size": "1000*-4016",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "1aacdc3de70a5217ef38d36f421e177d",
        "bound_box": "42,6292,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google account",
        "children": [
            372,
            373
        ],
        "focused": false,
        "bounds": [
            [
                42,
                6292
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 370,
        "temp_id": 371,
        "size": "1000*-4016",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "333c8aef9d2d8f54df46c20fd158e7e5",
        "bound_box": "42,6292,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                6344
            ],
            [
                916,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google account",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 371,
        "temp_id": 372,
        "size": "874*-4068",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Google account[enabled,,]",
        "view_str": "1850a24f0b38678b636305b72e192137",
        "bound_box": "42,6344,916,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                968,
                6344
            ],
            [
                1023,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.widget.Image",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 371,
        "temp_id": 373,
        "size": "55*-4068",
        "signature": "[class]android.widget.Image[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "8084260cfdf79c2c64e39058bd4490d5",
        "bound_box": "968,6344,1023,2276",
        "content_free_signature": "[class]android.widget.Image[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                6449
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 302,
        "temp_id": 374,
        "size": "1000*-4173",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "1b8d777b897133b175242f53ed4a7a08",
        "bound_box": "42,6449,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            376
        ],
        "focused": false,
        "bounds": [
            [
                42,
                6452
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": "2-0yZ-jtAcyGptQPofi-iA8__84",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 302,
        "temp_id": 375,
        "size": "1000*-4176",
        "signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__84[visible]False[text][enabled,,]",
        "view_str": "3d1f0484e4146d74d582e5d88377f3f5",
        "bound_box": "42,6452,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__84[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            377
        ],
        "focused": false,
        "bounds": [
            [
                42,
                6452
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 375,
        "temp_id": 376,
        "size": "1000*-4176",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "e0a299877010b054630a501c55a2b586",
        "bound_box": "42,6452,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "google.com search",
        "children": [
            378,
            379
        ],
        "focused": false,
        "bounds": [
            [
                42,
                6452
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 376,
        "temp_id": 377,
        "size": "1000*-4176",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "de3f1e6eef5900d9627febc79ff2fe63",
        "bound_box": "42,6452,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                6504
            ],
            [
                916,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "google.com search",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 377,
        "temp_id": 378,
        "size": "874*-4228",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]google.com search[enabled,,]",
        "view_str": "dfc5e6c2ca95c2737ae90ce8bd0becd4",
        "bound_box": "42,6504,916,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                968,
                6504
            ],
            [
                1023,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.widget.Image",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 377,
        "temp_id": 379,
        "size": "55*-4228",
        "signature": "[class]android.widget.Image[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "61ece082aae77147a56b749651896f3a",
        "bound_box": "968,6504,1023,2276",
        "content_free_signature": "[class]android.widget.Image[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                6609
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 302,
        "temp_id": 380,
        "size": "1000*-4333",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "1b8d777b897133b175242f53ed4a7a08",
        "bound_box": "42,6609,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            382
        ],
        "focused": false,
        "bounds": [
            [
                42,
                6612
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": "2-0yZ-jtAcyGptQPofi-iA8__86",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 302,
        "temp_id": 381,
        "size": "1000*-4336",
        "signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__86[visible]False[text][enabled,,]",
        "view_str": "98eff6b26857ba15ce500176f48198aa",
        "bound_box": "42,6612,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__86[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            383
        ],
        "focused": false,
        "bounds": [
            [
                42,
                6612
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 381,
        "temp_id": 382,
        "size": "1000*-4336",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "ed8a525a51bdfa5592100a684355a6e9",
        "bound_box": "42,6612,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google map",
        "children": [
            384,
            385
        ],
        "focused": false,
        "bounds": [
            [
                42,
                6612
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 382,
        "temp_id": 383,
        "size": "1000*-4336",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "14ffaa28f5447f5761c6d8fe6d09bf7f",
        "bound_box": "42,6612,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                6664
            ],
            [
                916,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google map",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 383,
        "temp_id": 384,
        "size": "874*-4388",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Google map[enabled,,]",
        "view_str": "36bfab7894cc4e29ac4376b813f5c998",
        "bound_box": "42,6664,916,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                968,
                6664
            ],
            [
                1023,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.widget.Image",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 383,
        "temp_id": 385,
        "size": "55*-4388",
        "signature": "[class]android.widget.Image[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "e50a420cce57d486be7c181064208ca4",
        "bound_box": "968,6664,1023,2276",
        "content_free_signature": "[class]android.widget.Image[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                6769
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 302,
        "temp_id": 386,
        "size": "1000*-4493",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "1b8d777b897133b175242f53ed4a7a08",
        "bound_box": "42,6769,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            388
        ],
        "focused": false,
        "bounds": [
            [
                42,
                6772
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": "2-0yZ-jtAcyGptQPofi-iA8__89",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 302,
        "temp_id": 387,
        "size": "1000*-4496",
        "signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__89[visible]False[text][enabled,,]",
        "view_str": "7f962e4ebb43b72d9bf7d9e938984a75",
        "bound_box": "42,6772,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__89[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            389
        ],
        "focused": false,
        "bounds": [
            [
                42,
                6772
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 387,
        "temp_id": 388,
        "size": "1000*-4496",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "042d9926f05ee32e1fb43c931c74f6ec",
        "bound_box": "42,6772,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google Mail",
        "children": [
            390,
            391
        ],
        "focused": false,
        "bounds": [
            [
                42,
                6772
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 388,
        "temp_id": 389,
        "size": "1000*-4496",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "cd9ab8cd5a5391628c37d31de4e808f5",
        "bound_box": "42,6772,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                6825
            ],
            [
                916,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google Mail",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 389,
        "temp_id": 390,
        "size": "874*-4549",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Google Mail[enabled,,]",
        "view_str": "7fea061e45e34d87004682d2a16a1b8a",
        "bound_box": "42,6825,916,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                968,
                6825
            ],
            [
                1023,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.widget.Image",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 389,
        "temp_id": 391,
        "size": "55*-4549",
        "signature": "[class]android.widget.Image[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "30dd4ed30f09c85d59f7043553222b28",
        "bound_box": "968,6825,1023,2276",
        "content_free_signature": "[class]android.widget.Image[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                -42,
                6930
            ],
            [
                1126,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 302,
        "temp_id": 392,
        "size": "1168*-4654",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "1b8d777b897133b175242f53ed4a7a08",
        "bound_box": "-42,6930,1126,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            394,
            396
        ],
        "focused": false,
        "bounds": [
            [
                0,
                6932
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 302,
        "temp_id": 393,
        "size": "1084*-4656",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "faecad1a71db4ad85580a054c89e7209",
        "bound_box": "0,6932,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            395
        ],
        "focused": false,
        "bounds": [
            [
                42,
                13678
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_137",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 393,
        "temp_id": 394,
        "size": "1000*-11402",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_137[visible]False[text][enabled,,]",
        "view_str": "b817f3295c5597c2e7e18e332d32ff37",
        "bound_box": "42,13678,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_137[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                6953
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_140",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 394,
        "temp_id": 395,
        "size": "1000*-4677",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_140[visible]False[text][enabled,,]",
        "view_str": "a9851b990855080eabd71050a3bf882a",
        "bound_box": "42,6953,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_140[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                882,
                6911
            ],
            [
                1063,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Feedback",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 393,
        "temp_id": 396,
        "size": "181*-4635",
        "signature": "[class]android.widget.Button[resource_id]None[visible]False[text]Feedback[enabled,,]",
        "view_str": "a598610a03d1bdd21cc99bc57c4530c5",
        "bound_box": "882,6911,1063,2276",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            398
        ],
        "focused": false,
        "bounds": [
            [
                0,
                7042
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 103,
        "temp_id": 397,
        "size": "1084*-4766",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "67049e768ef110aa9225cda8bf46cb44",
        "bound_box": "0,7042,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            399
        ],
        "focused": false,
        "bounds": [
            [
                0,
                7042
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 397,
        "temp_id": 398,
        "size": "1084*-4766",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "103594fa3687b9eb010a0cb55c42e6a8",
        "bound_box": "0,7042,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            400,
            410
        ],
        "focused": false,
        "bounds": [
            [
                0,
                7042
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 398,
        "temp_id": 399,
        "size": "1084*-4766",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "294a3a97a7aeea035b3f4a3ba19dbf29",
        "bound_box": "0,7042,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            401
        ],
        "focused": false,
        "bounds": [
            [
                0,
                7042
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 399,
        "temp_id": 400,
        "size": "1084*-4766",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "78957fc8d9d6bf28d42cd5753145ef6a",
        "bound_box": "0,7042,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 3,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            402,
            403,
            409
        ],
        "focused": false,
        "bounds": [
            [
                0,
                7042
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 400,
        "temp_id": 401,
        "size": "1084*-4766",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "d1d279c4989de55b621f270598adbeb2",
        "bound_box": "0,7042,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                7042
            ],
            [
                5,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Web results",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 401,
        "temp_id": 402,
        "size": "5*-4766",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Web results[enabled,,]",
        "view_str": "c8da96c4c07106792c13efb8f6ac6066",
        "bound_box": "0,7042,5,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google Blog https://blog.google › products › ge... Google Maps updates: Gemini arrives, Immersive View expands and more",
        "children": [
            404,
            408
        ],
        "focused": false,
        "bounds": [
            [
                0,
                7042
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 401,
        "temp_id": 403,
        "size": "1084*-4766",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "44c799870ddceb4be340e6670dcd371c",
        "bound_box": "0,7042,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            405
        ],
        "focused": false,
        "bounds": [
            [
                42,
                7082
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 403,
        "temp_id": 404,
        "size": "1000*-4806",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "14fc7afd7803359827765f00aca8214d",
        "bound_box": "42,7082,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            406,
            407
        ],
        "focused": false,
        "bounds": [
            [
                42,
                7082
            ],
            [
                937,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 404,
        "temp_id": 405,
        "size": "895*-4806",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "2f832e961eb8ab8151d44b648f7df66f",
        "bound_box": "42,7082,937,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                147,
                7084
            ],
            [
                658,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google Blog",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 405,
        "temp_id": 406,
        "size": "511*-4808",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Google Blog[enabled,,]",
        "view_str": "31d67341047fb3815771a5b578744a76",
        "bound_box": "147,7084,658,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                147,
                7140
            ],
            [
                658,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "https://blog.google › products › ge...",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 405,
        "temp_id": 407,
        "size": "511*-4864",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]https://blog.google › products › ge...[enabled,,]",
        "view_str": "68aa87b778a5e27210ce2340225153ba",
        "bound_box": "147,7140,658,2276",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                7210
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google Maps updates: Gemini arrives, Immersive View expands and more",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 403,
        "temp_id": 408,
        "size": "1000*-4934",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "d65c882daea8527e75ed186f714a0f7e",
        "bound_box": "42,7210,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                952,
                7042
            ],
            [
                1081,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "About this result",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 401,
        "temp_id": 409,
        "size": "129*-4766",
        "signature": "[class]android.widget.Button[resource_id]None[visible]False[text]About this result[enabled,,]",
        "view_str": "1664121feb337e00ea038619161786d9",
        "bound_box": "952,7042,1081,2276",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            411
        ],
        "focused": false,
        "bounds": [
            [
                0,
                7360
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 399,
        "temp_id": 410,
        "size": "1084*-5084",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "63bf2cd5a03b0f0b3405663df6b2874f",
        "bound_box": "0,7360,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                7365
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Oct 31, 2024 — From helping you explore even more with Immersive View to taking the stress out of your drive, here are updates on Google Maps you won't want to miss.",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 410,
        "temp_id": 411,
        "size": "1000*-5089",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "878c281d0b3766ccf7fdaeef4dec05b1",
        "bound_box": "42,7365,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                7575
            ],
            [
                5,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Twitter Results",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 103,
        "temp_id": 412,
        "size": "5*-5299",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Twitter Results[enabled,,]",
        "view_str": "3cde09d9bd34c2931ddd55351f057fbe",
        "bound_box": "0,7575,5,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            414
        ],
        "focused": false,
        "bounds": [
            [
                0,
                7575
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 103,
        "temp_id": 413,
        "size": "1084*-5299",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "67049e768ef110aa9225cda8bf46cb44",
        "bound_box": "0,7575,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            415,
            422
        ],
        "focused": false,
        "bounds": [
            [
                0,
                7575
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 413,
        "temp_id": 414,
        "size": "1084*-5299",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "ac20932b8aab54f5c24b10dd1c1529c4",
        "bound_box": "0,7575,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            416
        ],
        "focused": false,
        "bounds": [
            [
                0,
                7575
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 414,
        "temp_id": 415,
        "size": "1084*-5299",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "14377535e377fc74829bb389a08d7e9d",
        "bound_box": "0,7575,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            417,
            421
        ],
        "focused": false,
        "bounds": [
            [
                0,
                7575
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 415,
        "temp_id": 416,
        "size": "1084*-5299",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "c14915913789ae55d39336fe8457921b",
        "bound_box": "0,7575,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "X › Google Google",
        "children": [
            418,
            420
        ],
        "focused": false,
        "bounds": [
            [
                0,
                7575
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 416,
        "temp_id": 417,
        "size": "1084*-5299",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "4090d5f5cc4a915180c5ecb1748fc69a",
        "bound_box": "0,7575,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            419
        ],
        "focused": false,
        "bounds": [
            [
                42,
                7615
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 417,
        "temp_id": 418,
        "size": "1000*-5339",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "bf1bd2eff07cf022909e97947fb5c2aa",
        "bound_box": "42,7615,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                147,
                7625
            ],
            [
                294,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "X › Google",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 418,
        "temp_id": 419,
        "size": "147*-5349",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]X › Google[enabled,,]",
        "view_str": "730d3c6482391ace697f224c29e7b5a2",
        "bound_box": "147,7625,294,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                181,
                7720
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 417,
        "temp_id": 420,
        "size": "861*-5444",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Google[enabled,,]",
        "view_str": "473f198dd2970da5236746ae6e29396b",
        "bound_box": "181,7720,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                952,
                7575
            ],
            [
                1081,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "About this result",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 416,
        "temp_id": 421,
        "size": "129*-5299",
        "signature": "[class]android.widget.Button[resource_id]None[visible]False[text]About this result[enabled,,]",
        "view_str": "cf1824b6a44b6c942021738a366bafba",
        "bound_box": "952,7575,1081,2276",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            423
        ],
        "focused": false,
        "bounds": [
            [
                0,
                7827
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_113",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 414,
        "temp_id": 422,
        "size": "1084*-5551",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_113[visible]False[text][enabled,,]",
        "view_str": "afea94de0d7dc812251f7baadfe4b3b9",
        "bound_box": "0,7827,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_113[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            424
        ],
        "focused": false,
        "bounds": [
            [
                0,
                7827
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": true,
        "selected": false,
        "long_clickable": false,
        "parent": 422,
        "temp_id": 423,
        "size": "1084*-5551",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "9861c9540278d614ebb0f16f4efcd36e",
        "bound_box": "0,7827,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 6,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            425,
            437,
            450,
            463,
            478,
            491
        ],
        "focused": false,
        "bounds": [
            [
                42,
                7869
            ],
            [
                3480,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.widget.ListView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 423,
        "temp_id": 424,
        "size": "3438*-5593",
        "signature": "[class]android.widget.ListView[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "45fd1eae63062b407dd5185f8fc5e0a0",
        "bound_box": "42,7869,3480,2276",
        "content_free_signature": "[class]android.widget.ListView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            426
        ],
        "focused": false,
        "bounds": [
            [
                42,
                7869
            ],
            [
                640,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 424,
        "temp_id": 425,
        "size": "598*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "dc93076f0b2866a1d2657f5a37d254be",
        "bound_box": "42,7869,640,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            427
        ],
        "focused": false,
        "bounds": [
            [
                42,
                7869
            ],
            [
                640,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 425,
        "temp_id": 426,
        "size": "598*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "a6d493131d43e4eda305da913f9d7855",
        "bound_box": "42,7869,640,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            428
        ],
        "focused": false,
        "bounds": [
            [
                42,
                7869
            ],
            [
                640,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 426,
        "temp_id": 427,
        "size": "598*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "8c97ef5582654ce6deab22c9b2659fbe",
        "bound_box": "42,7869,640,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 3,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            429,
            430,
            436
        ],
        "focused": false,
        "bounds": [
            [
                42,
                7869
            ],
            [
                640,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 427,
        "temp_id": 428,
        "size": "598*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "a80771f1c56f8f6b35b928622cde9d58",
        "bound_box": "42,7869,640,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Floods cause catastrophic damage around the globe each year — but advance warnings can give people crucial time to take action before waters rise. Learn how we’re bringing our AI-powered flood forecasting to even more people ↓ goo.gle/3YMQ5Be",
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                7869
            ],
            [
                640,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 428,
        "temp_id": 429,
        "size": "598*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "5b047b669fca0df864c2e0211e1399a9",
        "bound_box": "42,7869,640,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            431
        ],
        "focused": false,
        "bounds": [
            [
                70,
                7898
            ],
            [
                606,
                2276
            ]
        ],
        "resource_id": "twitter_text_tsuid_2-0yZ-jtAcyGptQPofi-iA8_92",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 428,
        "temp_id": 430,
        "size": "536*-5622",
        "signature": "[class]android.view.View[resource_id]twitter_text_tsuid_2-0yZ-jtAcyGptQPofi-iA8_92[visible]False[text][enabled,,]",
        "view_str": "f100ca8370bbd54584a3d1cfbee8a974",
        "bound_box": "70,7898,606,2276",
        "content_free_signature": "[class]android.view.View[resource_id]twitter_text_tsuid_2-0yZ-jtAcyGptQPofi-iA8_92[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            432
        ],
        "focused": false,
        "bounds": [
            [
                70,
                7898
            ],
            [
                606,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 430,
        "temp_id": 431,
        "size": "536*-5622",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "e796304e50b077edd13831d807850f41",
        "bound_box": "70,7898,606,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            433,
            434
        ],
        "focused": false,
        "bounds": [
            [
                70,
                7898
            ],
            [
                606,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 431,
        "temp_id": 432,
        "size": "536*-5622",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "169382780580a2ee7a7dceaa28ac8663",
        "bound_box": "70,7898,606,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                70,
                7898
            ],
            [
                593,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Floods cause catastrophic damage around the globe each year — but advance warnings can give people crucial time to take action before waters rise. Learn how we’re bringing our AI-powered flood forecasting to even more people ↓ ",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 432,
        "temp_id": 433,
        "size": "523*-5622",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "305a071e79cda674964bb5731e668252",
        "bound_box": "70,7898,593,2276",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "goo.gle/3YMQ5Be",
        "children": [
            435
        ],
        "focused": false,
        "bounds": [
            [
                70,
                8276
            ],
            [
                378,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 432,
        "temp_id": 434,
        "size": "308*-6000",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "ce0eaa88603791af2a67e3df1927cb93",
        "bound_box": "70,8276,378,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                70,
                8276
            ],
            [
                378,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "goo.gle/3YMQ5Be",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 434,
        "temp_id": 435,
        "size": "308*-6000",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]goo.gle/3YMQ5Be[enabled,,]",
        "view_str": "f212faa1c179efbddce1338a73efb316",
        "bound_box": "70,8276,378,2276",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                70,
                8431
            ],
            [
                606,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "8 hours ago",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 428,
        "temp_id": 436,
        "size": "536*-6155",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]8 hours ago[enabled,,]",
        "view_str": "2da476ab272fdf705645bb34e6be23c5",
        "bound_box": "70,8431,606,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            438
        ],
        "focused": false,
        "bounds": [
            [
                666,
                7869
            ],
            [
                1265,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 424,
        "temp_id": 437,
        "size": "599*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "dc93076f0b2866a1d2657f5a37d254be",
        "bound_box": "666,7869,1265,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            439
        ],
        "focused": false,
        "bounds": [
            [
                666,
                7869
            ],
            [
                1265,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 437,
        "temp_id": 438,
        "size": "599*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "a6d493131d43e4eda305da913f9d7855",
        "bound_box": "666,7869,1265,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            440
        ],
        "focused": false,
        "bounds": [
            [
                666,
                7869
            ],
            [
                1265,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 438,
        "temp_id": 439,
        "size": "599*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "8c97ef5582654ce6deab22c9b2659fbe",
        "bound_box": "666,7869,1265,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 4,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            441,
            442,
            443,
            449
        ],
        "focused": false,
        "bounds": [
            [
                666,
                7869
            ],
            [
                1265,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 439,
        "temp_id": 440,
        "size": "599*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "a5d45b577c6fae2c3fba25e062ee80a0",
        "bound_box": "666,7869,1265,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "1856061214532465126?ref_src=twsrc%5Egoogle%7Ctwcamp%5Eserp%7Ctwgr%5Etweet",
        "children": [],
        "focused": false,
        "bounds": [
            [
                666,
                7869
            ],
            [
                1265,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 440,
        "temp_id": 441,
        "size": "599*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "5b047b669fca0df864c2e0211e1399a9",
        "bound_box": "666,7869,1265,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Vets who own small businesses can join our #NationalVeteransSmallBusinessWeek Virtual Summit on Nov 13, hosted by #GrowWithGoogle and @BlueStarFamily to learn how our AI tools can help improve efficiency, customer service and more → g.co/grow/NVSBW",
        "children": [],
        "focused": false,
        "bounds": [
            [
                666,
                7869
            ],
            [
                1265,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 440,
        "temp_id": 442,
        "size": "599*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "5b047b669fca0df864c2e0211e1399a9",
        "bound_box": "666,7869,1265,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            444
        ],
        "focused": false,
        "bounds": [
            [
                698,
                8221
            ],
            [
                1233,
                2276
            ]
        ],
        "resource_id": "twitter_text_tsuid_2-0yZ-jtAcyGptQPofi-iA8_95",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 440,
        "temp_id": 443,
        "size": "535*-5945",
        "signature": "[class]android.view.View[resource_id]twitter_text_tsuid_2-0yZ-jtAcyGptQPofi-iA8_95[visible]False[text][enabled,,]",
        "view_str": "7fa313c1c57487282ac8c5c4ab10870b",
        "bound_box": "698,8221,1233,2276",
        "content_free_signature": "[class]android.view.View[resource_id]twitter_text_tsuid_2-0yZ-jtAcyGptQPofi-iA8_95[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            445
        ],
        "focused": false,
        "bounds": [
            [
                698,
                8221
            ],
            [
                1233,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 443,
        "temp_id": 444,
        "size": "535*-5945",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "d4044a7ed63d96bfa19e0bf7424ecb07",
        "bound_box": "698,8221,1233,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            446,
            447
        ],
        "focused": false,
        "bounds": [
            [
                698,
                8221
            ],
            [
                1233,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 444,
        "temp_id": 445,
        "size": "535*-5945",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "059ca819c9f3a62d12d39cf5038c6c80",
        "bound_box": "698,8221,1233,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                698,
                8221
            ],
            [
                1330,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Vets who own small businesses can join our #NationalVeteransSmallBusinessWeek Virtual Summit on Nov 13, hosted by #GrowWithGoogle and @BlueStarFamily to learn how our AI tools can help improve efficiency, customer service and more → ",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 445,
        "temp_id": 446,
        "size": "632*-5945",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "0149c46b475a329837d91abae0daaf46",
        "bound_box": "698,8221,1330,2276",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "g.co/grow/NVSBW",
        "children": [
            448
        ],
        "focused": false,
        "bounds": [
            [
                698,
                8646
            ],
            [
                1002,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 445,
        "temp_id": 447,
        "size": "304*-6370",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "55da5fa7c2d6c458a8b2c1b33e771909",
        "bound_box": "698,8646,1002,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                698,
                8646
            ],
            [
                1002,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "g.co/grow/NVSBW",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 447,
        "temp_id": 448,
        "size": "304*-6370",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]g.co/grow/NVSBW[enabled,,]",
        "view_str": "c31d5cc78c11057c08b7979c3c8091b5",
        "bound_box": "698,8646,1002,2276",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                698,
                8431
            ],
            [
                1233,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "10 hours ago",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 440,
        "temp_id": 449,
        "size": "535*-6155",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]10 hours ago[enabled,,]",
        "view_str": "a295d70098848636058acbe44c33c77b",
        "bound_box": "698,8431,1233,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            451
        ],
        "focused": false,
        "bounds": [
            [
                1294,
                7869
            ],
            [
                1892,
                2276
            ]
        ],
        "resource_id": "tsuid_2-0yZ-jtAcyGptQPofi-iA8_114",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 424,
        "temp_id": 450,
        "size": "598*-5593",
        "signature": "[class]android.view.View[resource_id]tsuid_2-0yZ-jtAcyGptQPofi-iA8_114[visible]False[text][enabled,,]",
        "view_str": "18b18ba290b236680a0eb0f6ebf98e25",
        "bound_box": "1294,7869,1892,2276",
        "content_free_signature": "[class]android.view.View[resource_id]tsuid_2-0yZ-jtAcyGptQPofi-iA8_114[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            452
        ],
        "focused": false,
        "bounds": [
            [
                1294,
                7869
            ],
            [
                1892,
                2276
            ]
        ],
        "resource_id": "2-0yZ-jtAcyGptQPofi-iA8__58",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 450,
        "temp_id": 451,
        "size": "598*-5593",
        "signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__58[visible]False[text][enabled,,]",
        "view_str": "28db653c6f796d7f39214e2ea9d2d18b",
        "bound_box": "1294,7869,1892,2276",
        "content_free_signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__58[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            453
        ],
        "focused": false,
        "bounds": [
            [
                1294,
                7869
            ],
            [
                1892,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 451,
        "temp_id": 452,
        "size": "598*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "33e16cb7008f4a0fa432a74055fa69ff",
        "bound_box": "1294,7869,1892,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            454
        ],
        "focused": false,
        "bounds": [
            [
                1294,
                7869
            ],
            [
                1892,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 452,
        "temp_id": 453,
        "size": "598*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "8a7f061329eb95368eb05a01e995716f",
        "bound_box": "1294,7869,1892,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 3,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            455,
            456,
            462
        ],
        "focused": false,
        "bounds": [
            [
                1294,
                7869
            ],
            [
                1892,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 453,
        "temp_id": 454,
        "size": "598*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "e8d7dc9cd0c5cf667ff909ab02f5af81",
        "bound_box": "1294,7869,1892,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "This #VeteransDay, we’re honoring the contributions of veterans and their families, as well as highlighting programs Googlers launched this year to empower vets as they transition into life as civilians. Here’s how ↓ goo.gle/4fm4xYb",
        "children": [],
        "focused": false,
        "bounds": [
            [
                1294,
                7869
            ],
            [
                1892,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 454,
        "temp_id": 455,
        "size": "598*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "184f8637f4242ec69cc99bef67a4528c",
        "bound_box": "1294,7869,1892,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            457
        ],
        "focused": false,
        "bounds": [
            [
                1325,
                7898
            ],
            [
                1861,
                2276
            ]
        ],
        "resource_id": "twitter_text_tsuid_2-0yZ-jtAcyGptQPofi-iA8_98",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 454,
        "temp_id": 456,
        "size": "536*-5622",
        "signature": "[class]android.view.View[resource_id]twitter_text_tsuid_2-0yZ-jtAcyGptQPofi-iA8_98[visible]False[text][enabled,,]",
        "view_str": "4722c17ad359a09a0d395e64cd0e10ec",
        "bound_box": "1325,7898,1861,2276",
        "content_free_signature": "[class]android.view.View[resource_id]twitter_text_tsuid_2-0yZ-jtAcyGptQPofi-iA8_98[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            458
        ],
        "focused": false,
        "bounds": [
            [
                1325,
                7898
            ],
            [
                1861,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 456,
        "temp_id": 457,
        "size": "536*-5622",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "3311c455df478d4ba0bb11da4e637aa7",
        "bound_box": "1325,7898,1861,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            459,
            460
        ],
        "focused": false,
        "bounds": [
            [
                1325,
                7898
            ],
            [
                1861,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 457,
        "temp_id": 458,
        "size": "536*-5622",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "d5a850c976230ad9f5c3012ea60864fa",
        "bound_box": "1325,7898,1861,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1325,
                7898
            ],
            [
                1858,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "This #VeteransDay, we’re honoring the contributions of veterans and their families, as well as highlighting programs Googlers launched this year to empower vets as they transition into life as civilians. Here’s how ↓ ",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 458,
        "temp_id": 459,
        "size": "533*-5622",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "4109b2b8a47d59946c10e9bf6dddd759",
        "bound_box": "1325,7898,1858,2276",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "goo.gle/4fm4xYb",
        "children": [
            461
        ],
        "focused": false,
        "bounds": [
            [
                1325,
                8229
            ],
            [
                1611,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 458,
        "temp_id": 460,
        "size": "286*-5953",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "0d9f018221120b82c9b3e38fa4a3c76d",
        "bound_box": "1325,8229,1611,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1325,
                8229
            ],
            [
                1611,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "goo.gle/4fm4xYb",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 460,
        "temp_id": 461,
        "size": "286*-5953",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]goo.gle/4fm4xYb[enabled,,]",
        "view_str": "d7cdc7da69a2bc222f10df8376639616",
        "bound_box": "1325,8229,1611,2276",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1325,
                8431
            ],
            [
                1861,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "15 hours ago",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 454,
        "temp_id": 462,
        "size": "536*-6155",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]15 hours ago[enabled,,]",
        "view_str": "31278066a1502c9674df5c7db7ff107a",
        "bound_box": "1325,8431,1861,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            464
        ],
        "focused": false,
        "bounds": [
            [
                1918,
                7869
            ],
            [
                2517,
                2276
            ]
        ],
        "resource_id": "tsuid_2-0yZ-jtAcyGptQPofi-iA8_116",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 424,
        "temp_id": 463,
        "size": "599*-5593",
        "signature": "[class]android.view.View[resource_id]tsuid_2-0yZ-jtAcyGptQPofi-iA8_116[visible]False[text][enabled,,]",
        "view_str": "005f1d5e9f6baa1051dca8adf4485760",
        "bound_box": "1918,7869,2517,2276",
        "content_free_signature": "[class]android.view.View[resource_id]tsuid_2-0yZ-jtAcyGptQPofi-iA8_116[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            465
        ],
        "focused": false,
        "bounds": [
            [
                1918,
                7869
            ],
            [
                2517,
                2276
            ]
        ],
        "resource_id": "2-0yZ-jtAcyGptQPofi-iA8__60",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 463,
        "temp_id": 464,
        "size": "599*-5593",
        "signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__60[visible]False[text][enabled,,]",
        "view_str": "132ebc8ef89c85f86c1f1c0decb3adc1",
        "bound_box": "1918,7869,2517,2276",
        "content_free_signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__60[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            466
        ],
        "focused": false,
        "bounds": [
            [
                1918,
                7869
            ],
            [
                2517,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 464,
        "temp_id": 465,
        "size": "599*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "a34bb2e135916bcf7ed16db3e80d8911",
        "bound_box": "1918,7869,2517,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            467
        ],
        "focused": false,
        "bounds": [
            [
                1918,
                7869
            ],
            [
                2517,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 465,
        "temp_id": 466,
        "size": "599*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "7d3a9db62d8f468a06ac3fc8df52f255",
        "bound_box": "1918,7869,2517,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 4,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            468,
            469,
            470,
            477
        ],
        "focused": false,
        "bounds": [
            [
                1918,
                7869
            ],
            [
                2517,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 466,
        "temp_id": 467,
        "size": "599*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "c570027344087c722513dd7ca1ca2e9b",
        "bound_box": "1918,7869,2517,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "1854646590113304589?ref_src=twsrc%5Egoogle%7Ctwcamp%5Eserp%7Ctwgr%5Etweet",
        "children": [],
        "focused": false,
        "bounds": [
            [
                1918,
                7869
            ],
            [
                2517,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 467,
        "temp_id": 468,
        "size": "599*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "702fc99cbfa09b4fc97f8ffd281d42c0",
        "bound_box": "1918,7869,2517,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Get ready for the GRAMMYs nominations, streaming live on @YouTube on Friday, 11/8 at 11 a.m. ET → yt.be/grammys Who do you think should be nominated?",
        "children": [],
        "focused": false,
        "bounds": [
            [
                1918,
                7869
            ],
            [
                2517,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 467,
        "temp_id": 469,
        "size": "599*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "702fc99cbfa09b4fc97f8ffd281d42c0",
        "bound_box": "1918,7869,2517,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            471
        ],
        "focused": false,
        "bounds": [
            [
                1953,
                8221
            ],
            [
                2488,
                2276
            ]
        ],
        "resource_id": "twitter_text_tsuid_2-0yZ-jtAcyGptQPofi-iA8_100",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 467,
        "temp_id": 470,
        "size": "535*-5945",
        "signature": "[class]android.view.View[resource_id]twitter_text_tsuid_2-0yZ-jtAcyGptQPofi-iA8_100[visible]False[text][enabled,,]",
        "view_str": "3e2b8353affe60977b65d3b71febec9f",
        "bound_box": "1953,8221,2488,2276",
        "content_free_signature": "[class]android.view.View[resource_id]twitter_text_tsuid_2-0yZ-jtAcyGptQPofi-iA8_100[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            472
        ],
        "focused": false,
        "bounds": [
            [
                1953,
                8221
            ],
            [
                2488,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 470,
        "temp_id": 471,
        "size": "535*-5945",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "8deb8dae19dd27556fa2971d38ebbbcb",
        "bound_box": "1953,8221,2488,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 3,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            473,
            474,
            476
        ],
        "focused": false,
        "bounds": [
            [
                1953,
                8221
            ],
            [
                2488,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 471,
        "temp_id": 472,
        "size": "535*-5945",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "409e77cd3d8c78c7577619813a3b8ef2",
        "bound_box": "1953,8221,2488,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1953,
                8221
            ],
            [
                2457,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Get ready for the GRAMMYs nominations, streaming live on @YouTube on Friday, 11/8 at 11 a.m. ET → ",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 472,
        "temp_id": 473,
        "size": "504*-5945",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "773752c4c46a6ab9661e9c708a366013",
        "bound_box": "1953,8221,2457,2276",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "yt.be/grammys",
        "children": [
            475
        ],
        "focused": false,
        "bounds": [
            [
                2123,
                8363
            ],
            [
                2373,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 472,
        "temp_id": 474,
        "size": "250*-6087",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "761492b09175ff10397ac994c4a3aaa6",
        "bound_box": "2123,8363,2373,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                2123,
                8363
            ],
            [
                2373,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "yt.be/grammys",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 474,
        "temp_id": 475,
        "size": "250*-6087",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]yt.be/grammys[enabled,,]",
        "view_str": "b0394ec5c1dc7f81b446903a01bae082",
        "bound_box": "2123,8363,2373,2276",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1953,
                8363
            ],
            [
                2415,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "\nWho do you think should be nominated?",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 472,
        "temp_id": 476,
        "size": "462*-6087",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]\nWho do you think should be nominated?[enabled,,]",
        "view_str": "d782d747ae0f6207c11b924b0fc4cad1",
        "bound_box": "1953,8363,2415,2276",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1953,
                8431
            ],
            [
                2488,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "4 days ago",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 467,
        "temp_id": 477,
        "size": "535*-6155",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]4 days ago[enabled,,]",
        "view_str": "6def812c651a8b30bbd8454d248c20df",
        "bound_box": "1953,8431,2488,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            479
        ],
        "focused": false,
        "bounds": [
            [
                2546,
                7869
            ],
            [
                3144,
                2276
            ]
        ],
        "resource_id": "tsuid_2-0yZ-jtAcyGptQPofi-iA8_119",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 424,
        "temp_id": 478,
        "size": "598*-5593",
        "signature": "[class]android.view.View[resource_id]tsuid_2-0yZ-jtAcyGptQPofi-iA8_119[visible]False[text][enabled,,]",
        "view_str": "2bc22f888b6df66506dfd9c19d1a55de",
        "bound_box": "2546,7869,3144,2276",
        "content_free_signature": "[class]android.view.View[resource_id]tsuid_2-0yZ-jtAcyGptQPofi-iA8_119[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            480
        ],
        "focused": false,
        "bounds": [
            [
                2546,
                7869
            ],
            [
                3144,
                2276
            ]
        ],
        "resource_id": "2-0yZ-jtAcyGptQPofi-iA8__62",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 478,
        "temp_id": 479,
        "size": "598*-5593",
        "signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__62[visible]False[text][enabled,,]",
        "view_str": "fd44e458b18325c04e415631bedd0315",
        "bound_box": "2546,7869,3144,2276",
        "content_free_signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__62[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            481
        ],
        "focused": false,
        "bounds": [
            [
                2546,
                7869
            ],
            [
                3144,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 479,
        "temp_id": 480,
        "size": "598*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "830e4ae9a30a45db830b942f9dad5a49",
        "bound_box": "2546,7869,3144,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            482
        ],
        "focused": false,
        "bounds": [
            [
                2546,
                7869
            ],
            [
                3144,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 480,
        "temp_id": 481,
        "size": "598*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "80ccf4de067251ab6f14c74d5dcb449d",
        "bound_box": "2546,7869,3144,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 3,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            483,
            484,
            490
        ],
        "focused": false,
        "bounds": [
            [
                2546,
                7869
            ],
            [
                3144,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 481,
        "temp_id": 482,
        "size": "598*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "d3e0a769ed050488db29cfe5ebbfcfa5",
        "bound_box": "2546,7869,3144,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Catch up on our latest AI updates from October 🛍️ Find products you love with new Shopping features 🔎 New ways to search, like video in Lens 🚘 An even more helpful Maps And more ↓ goo.gle/3YyUzva",
        "children": [],
        "focused": false,
        "bounds": [
            [
                2546,
                7869
            ],
            [
                3144,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 482,
        "temp_id": 483,
        "size": "598*-5593",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "a1989ebe281123b4fa0281649a63d67e",
        "bound_box": "2546,7869,3144,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            485
        ],
        "focused": false,
        "bounds": [
            [
                2577,
                7898
            ],
            [
                3113,
                2276
            ]
        ],
        "resource_id": "twitter_text_tsuid_2-0yZ-jtAcyGptQPofi-iA8_96",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 482,
        "temp_id": 484,
        "size": "536*-5622",
        "signature": "[class]android.view.View[resource_id]twitter_text_tsuid_2-0yZ-jtAcyGptQPofi-iA8_96[visible]False[text][enabled,,]",
        "view_str": "e5b71b6abe46d070716c884985644ee0",
        "bound_box": "2577,7898,3113,2276",
        "content_free_signature": "[class]android.view.View[resource_id]twitter_text_tsuid_2-0yZ-jtAcyGptQPofi-iA8_96[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            486
        ],
        "focused": false,
        "bounds": [
            [
                2577,
                7898
            ],
            [
                3113,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 484,
        "temp_id": 485,
        "size": "536*-5622",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "a410963c1b4aaab9fb2e81d0003429bb",
        "bound_box": "2577,7898,3113,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            487,
            488
        ],
        "focused": false,
        "bounds": [
            [
                2577,
                7898
            ],
            [
                3113,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 485,
        "temp_id": 486,
        "size": "536*-5622",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "22bf025512c41d4365095817ca64f5f6",
        "bound_box": "2577,7898,3113,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                2577,
                7898
            ],
            [
                3089,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Catch up on our latest AI updates from October\n🛍️ Find products you love with new Shopping features\n🔎 New ways to search, like video in Lens\n🚘 An even more helpful Maps\nAnd more ↓\n",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 486,
        "temp_id": 487,
        "size": "512*-5622",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "b8968296493f3ec98f588438a9f714f4",
        "bound_box": "2577,7898,3089,2276",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "goo.gle/3YyUzva",
        "children": [
            489
        ],
        "focused": false,
        "bounds": [
            [
                2577,
                8276
            ],
            [
                2856,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 486,
        "temp_id": 488,
        "size": "279*-6000",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "40e623d2e8070a6f4e8e52f36b5964de",
        "bound_box": "2577,8276,2856,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                2577,
                8276
            ],
            [
                2856,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "goo.gle/3YyUzva",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 488,
        "temp_id": 489,
        "size": "279*-6000",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]goo.gle/3YyUzva[enabled,,]",
        "view_str": "4492a1461014e250175d82cb71b63843",
        "bound_box": "2577,8276,2856,2276",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                2577,
                8431
            ],
            [
                3113,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Nov 1, 2024",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 482,
        "temp_id": 490,
        "size": "536*-6155",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Nov 1, 2024[enabled,,]",
        "view_str": "dd2e7003a1821637a842a48b1bc6dda4",
        "bound_box": "2577,8431,3113,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            492
        ],
        "focused": false,
        "bounds": [
            [
                3173,
                7869
            ],
            [
                3507,
                2276
            ]
        ],
        "resource_id": "tsuid_2-0yZ-jtAcyGptQPofi-iA8_121",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 424,
        "temp_id": 491,
        "size": "334*-5593",
        "signature": "[class]android.view.View[resource_id]tsuid_2-0yZ-jtAcyGptQPofi-iA8_121[visible]False[text][enabled,,]",
        "view_str": "558949a2263162a5780fffc602bd1c03",
        "bound_box": "3173,7869,3507,2276",
        "content_free_signature": "[class]android.view.View[resource_id]tsuid_2-0yZ-jtAcyGptQPofi-iA8_121[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            493
        ],
        "focused": false,
        "bounds": [
            [
                3257,
                8095
            ],
            [
                3423,
                2276
            ]
        ],
        "resource_id": "2-0yZ-jtAcyGptQPofi-iA8__51",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 491,
        "temp_id": 492,
        "size": "166*-5819",
        "signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__51[visible]False[text][enabled,,]",
        "view_str": "e5d538e89405bd0bb58d3c5174a14949",
        "bound_box": "3257,8095,3423,2276",
        "content_free_signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__51[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "View on X",
        "children": [
            494
        ],
        "focused": false,
        "bounds": [
            [
                3257,
                8095
            ],
            [
                3423,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 492,
        "temp_id": 493,
        "size": "166*-5819",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "8c0e00efcbcda2f86af5792d89dcddeb",
        "bound_box": "3257,8095,3423,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            495,
            497
        ],
        "focused": false,
        "bounds": [
            [
                3257,
                8095
            ],
            [
                3423,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 493,
        "temp_id": 494,
        "size": "166*-5819",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "ec747b32820768d1910dc4fc13bcf176",
        "bound_box": "3257,8095,3423,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            496
        ],
        "focused": false,
        "bounds": [
            [
                3281,
                8095
            ],
            [
                3399,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 494,
        "temp_id": 495,
        "size": "118*-5819",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "b940198a5a55952309a537495e011de3",
        "bound_box": "3281,8095,3399,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                3312,
                8127
            ],
            [
                3367,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.widget.Image",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 495,
        "temp_id": 496,
        "size": "55*-5851",
        "signature": "[class]android.widget.Image[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "59f8a0fdb3477db8b8c63480da8396c7",
        "bound_box": "3312,8127,3367,2276",
        "content_free_signature": "[class]android.widget.Image[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                3257,
                8226
            ],
            [
                3423,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "View on X",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 494,
        "temp_id": 497,
        "size": "166*-5950",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]View on X[enabled,,]",
        "view_str": "1758b0bf92940cd6b0773fc95816cf78",
        "bound_box": "3257,8226,3423,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            499
        ],
        "focused": false,
        "bounds": [
            [
                0,
                8568
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 103,
        "temp_id": 498,
        "size": "1084*-6292",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "67049e768ef110aa9225cda8bf46cb44",
        "bound_box": "0,8568,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            500
        ],
        "focused": false,
        "bounds": [
            [
                0,
                8568
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 498,
        "temp_id": 499,
        "size": "1084*-6292",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "103594fa3687b9eb010a0cb55c42e6a8",
        "bound_box": "0,8568,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            501,
            511
        ],
        "focused": false,
        "bounds": [
            [
                0,
                8568
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 499,
        "temp_id": 500,
        "size": "1084*-6292",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "294a3a97a7aeea035b3f4a3ba19dbf29",
        "bound_box": "0,8568,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            502
        ],
        "focused": false,
        "bounds": [
            [
                0,
                8568
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 500,
        "temp_id": 501,
        "size": "1084*-6292",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "78957fc8d9d6bf28d42cd5753145ef6a",
        "bound_box": "0,8568,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 3,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            503,
            504,
            510
        ],
        "focused": false,
        "bounds": [
            [
                0,
                8568
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 501,
        "temp_id": 502,
        "size": "1084*-6292",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "d1d279c4989de55b621f270598adbeb2",
        "bound_box": "0,8568,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                8568
            ],
            [
                5,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Web results",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 502,
        "temp_id": 503,
        "size": "5*-6292",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Web results[enabled,,]",
        "view_str": "c8da96c4c07106792c13efb8f6ac6066",
        "bound_box": "0,8568,5,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "About Google https://about.google Google - About Google, Our Culture & Company News",
        "children": [
            505,
            509
        ],
        "focused": false,
        "bounds": [
            [
                0,
                8568
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 502,
        "temp_id": 504,
        "size": "1084*-6292",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "50224b70c5a03af2cbaecd8fb90914ef",
        "bound_box": "0,8568,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            506
        ],
        "focused": false,
        "bounds": [
            [
                42,
                8607
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 504,
        "temp_id": 505,
        "size": "1000*-6331",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "14fc7afd7803359827765f00aca8214d",
        "bound_box": "42,8607,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            507,
            508
        ],
        "focused": false,
        "bounds": [
            [
                42,
                8607
            ],
            [
                937,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 505,
        "temp_id": 506,
        "size": "895*-6331",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "c8764023b787915ca4c1702011cbdc2d",
        "bound_box": "42,8607,937,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                147,
                8610
            ],
            [
                441,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "About Google",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 506,
        "temp_id": 507,
        "size": "294*-6334",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]About Google[enabled,,]",
        "view_str": "06acb0c5f002e7d282f527b5bf8c4382",
        "bound_box": "147,8610,441,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                147,
                8667
            ],
            [
                441,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "https://about.google",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 506,
        "temp_id": 508,
        "size": "294*-6391",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]https://about.google[enabled,,]",
        "view_str": "762bf5b4115a5441f8e1f434e85d6dfa",
        "bound_box": "147,8667,441,2276",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                8736
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google - About Google, Our Culture & Company News",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 504,
        "temp_id": 509,
        "size": "1000*-6460",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Google - About Google, Our Culture & Company News[enabled,,]",
        "view_str": "9394647762910ff6f4e1d3ed204128ca",
        "bound_box": "42,8736,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                952,
                8568
            ],
            [
                1081,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "About this result",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 502,
        "temp_id": 510,
        "size": "129*-6292",
        "signature": "[class]android.widget.Button[resource_id]None[visible]False[text]About this result[enabled,,]",
        "view_str": "1664121feb337e00ea038619161786d9",
        "bound_box": "952,8568,1081,2276",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            512
        ],
        "focused": false,
        "bounds": [
            [
                0,
                8885
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 500,
        "temp_id": 511,
        "size": "1084*-6609",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "63bf2cd5a03b0f0b3405663df6b2874f",
        "bound_box": "0,8885,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                8890
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Stay up to date with Google company news and products. Discover stories about our culture, philosophy, and how Google technology is impacting others.",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 511,
        "temp_id": 512,
        "size": "1000*-6614",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "878c281d0b3766ccf7fdaeef4dec05b1",
        "bound_box": "42,8890,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            514
        ],
        "focused": false,
        "bounds": [
            [
                0,
                9100
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 103,
        "temp_id": 513,
        "size": "1084*-6824",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "67049e768ef110aa9225cda8bf46cb44",
        "bound_box": "0,9100,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            515
        ],
        "focused": false,
        "bounds": [
            [
                0,
                9100
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 513,
        "temp_id": 514,
        "size": "1084*-6824",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "103594fa3687b9eb010a0cb55c42e6a8",
        "bound_box": "0,9100,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 3,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            516,
            525,
            527
        ],
        "focused": false,
        "bounds": [
            [
                0,
                9100
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 514,
        "temp_id": 515,
        "size": "1084*-6824",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "af4a96a71350767ffda65ff752b99edf",
        "bound_box": "0,9100,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            517
        ],
        "focused": false,
        "bounds": [
            [
                0,
                9100
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 515,
        "temp_id": 516,
        "size": "1084*-6824",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "78957fc8d9d6bf28d42cd5753145ef6a",
        "bound_box": "0,9100,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            518,
            524
        ],
        "focused": false,
        "bounds": [
            [
                0,
                9100
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 516,
        "temp_id": 517,
        "size": "1084*-6824",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "9059e8fff283cdedad5a4073a983c285",
        "bound_box": "0,9100,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Wikipedia https://en.wikipedia.org › wiki › G... Google",
        "children": [
            519,
            523
        ],
        "focused": false,
        "bounds": [
            [
                0,
                9100
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 517,
        "temp_id": 518,
        "size": "1084*-6824",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "0d81c960d94864d0cfdcc5e0142008a6",
        "bound_box": "0,9100,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            520
        ],
        "focused": false,
        "bounds": [
            [
                42,
                9140
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 518,
        "temp_id": 519,
        "size": "1000*-6864",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "14fc7afd7803359827765f00aca8214d",
        "bound_box": "42,9140,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            521,
            522
        ],
        "focused": false,
        "bounds": [
            [
                42,
                9140
            ],
            [
                937,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 519,
        "temp_id": 520,
        "size": "895*-6864",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "98a7ab7443d9d7bd68f4d82c2b1037f8",
        "bound_box": "42,9140,937,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                147,
                9142
            ],
            [
                640,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Wikipedia",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 520,
        "temp_id": 521,
        "size": "493*-6866",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Wikipedia[enabled,,]",
        "view_str": "05fb36c5876eef51a1852716c6e35781",
        "bound_box": "147,9142,640,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                147,
                9198
            ],
            [
                640,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "https://en.wikipedia.org › wiki › G...",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 520,
        "temp_id": 522,
        "size": "493*-6922",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]https://en.wikipedia.org › wiki › G...[enabled,,]",
        "view_str": "f20912635ccd4ce1364d2365be4fc7e4",
        "bound_box": "147,9198,640,2276",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                9268
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 518,
        "temp_id": 523,
        "size": "1000*-6992",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Google[enabled,,]",
        "view_str": "69321ac291960a8357cad1338c8592e8",
        "bound_box": "42,9268,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                952,
                9100
            ],
            [
                1081,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "About this result",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 517,
        "temp_id": 524,
        "size": "129*-6824",
        "signature": "[class]android.widget.Button[resource_id]None[visible]False[text]About this result[enabled,,]",
        "view_str": "1664121feb337e00ea038619161786d9",
        "bound_box": "952,9100,1081,2276",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            526
        ],
        "focused": false,
        "bounds": [
            [
                0,
                9352
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 515,
        "temp_id": 525,
        "size": "1084*-7076",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "63bf2cd5a03b0f0b3405663df6b2874f",
        "bound_box": "0,9352,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                9355
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google LLC is an American-based multinational corporation and technology company focusing on online advertising, search engine technology, cloud computing, ...",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 525,
        "temp_id": 526,
        "size": "1000*-7079",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "878c281d0b3766ccf7fdaeef4dec05b1",
        "bound_box": "42,9355,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            528
        ],
        "focused": false,
        "bounds": [
            [
                0,
                9528
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 515,
        "temp_id": 527,
        "size": "1084*-7252",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "78957fc8d9d6bf28d42cd5753145ef6a",
        "bound_box": "0,9528,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            529
        ],
        "focused": false,
        "bounds": [
            [
                0,
                9544
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 527,
        "temp_id": 528,
        "size": "1084*-7268",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "115268acf822c3866e5eb7f133f34992",
        "bound_box": "0,9544,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            530
        ],
        "focused": false,
        "bounds": [
            [
                0,
                9544
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": true,
        "selected": false,
        "long_clickable": false,
        "parent": 528,
        "temp_id": 529,
        "size": "1084*-7268",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "571457d2e2dc2d5c0c79b5abc5f729af",
        "bound_box": "0,9544,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 7,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            531,
            533,
            535,
            537,
            539,
            541,
            543
        ],
        "focused": false,
        "bounds": [
            [
                0,
                9544
            ],
            [
                2336,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 529,
        "temp_id": 530,
        "size": "2336*-7268",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "fe2d825f68a3639c3f6b85583bce2e62",
        "bound_box": "0,9544,2336,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "History",
        "children": [
            532
        ],
        "focused": false,
        "bounds": [
            [
                42,
                9544
            ],
            [
                231,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 530,
        "temp_id": 531,
        "size": "189*-7268",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "ed97a9b5300e958a1297596f5e010b1f",
        "bound_box": "42,9544,231,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                9544
            ],
            [
                231,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "History",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 531,
        "temp_id": 532,
        "size": "189*-7268",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]History[enabled,,]",
        "view_str": "584380ddaa8abf598962a4b3e9ebfd83",
        "bound_box": "42,9544,231,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google Chrome",
        "children": [
            534
        ],
        "focused": false,
        "bounds": [
            [
                225,
                9544
            ],
            [
                569,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 530,
        "temp_id": 533,
        "size": "344*-7268",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "1d4d6e2e9960d7a1a8221db15e818513",
        "bound_box": "225,9544,569,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                241,
                9544
            ],
            [
                569,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google Chrome",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 533,
        "temp_id": 534,
        "size": "328*-7268",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Google Chrome[enabled,,]",
        "view_str": "3d6f8a1e8bc6c14bffb50f6ca39dc2a2",
        "bound_box": "241,9544,569,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google Pixel",
        "children": [
            536
        ],
        "focused": false,
        "bounds": [
            [
                567,
                9544
            ],
            [
                858,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 530,
        "temp_id": 535,
        "size": "291*-7268",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "54d8e4299ea31019ff70aa7ea3be0188",
        "bound_box": "567,9544,858,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                582,
                9544
            ],
            [
                858,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google Pixel",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 535,
        "temp_id": 536,
        "size": "276*-7268",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Google Pixel[enabled,,]",
        "view_str": "995ea096e27c73dd4c2c2b76c4ff35e8",
        "bound_box": "582,9544,858,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google Nest",
        "children": [
            538
        ],
        "focused": false,
        "bounds": [
            [
                855,
                9544
            ],
            [
                1147,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 530,
        "temp_id": 537,
        "size": "292*-7268",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "9702aa7c97c418e12455c422932a4e42",
        "bound_box": "855,9544,1147,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                871,
                9544
            ],
            [
                1147,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google Nest",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 537,
        "temp_id": 538,
        "size": "276*-7268",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Google Nest[enabled,,]",
        "view_str": "cbd8f6f17c28103a5cf3840c94c67b29",
        "bound_box": "871,9544,1147,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google (disambiguation)",
        "children": [
            540
        ],
        "focused": false,
        "bounds": [
            [
                1141,
                9544
            ],
            [
                1635,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 530,
        "temp_id": 539,
        "size": "494*-7268",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "f7fb5ffe2c43923167ffad078f01a07e",
        "bound_box": "1141,9544,1635,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1157,
                9544
            ],
            [
                1635,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google (disambiguation)",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 539,
        "temp_id": 540,
        "size": "478*-7268",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Google (disambiguation)[enabled,,]",
        "view_str": "f5c8ff9b99759207efe5b03845fc4bd3",
        "bound_box": "1157,9544,1635,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google DeepMind",
        "children": [
            542
        ],
        "focused": false,
        "bounds": [
            [
                1632,
                9544
            ],
            [
                2013,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 530,
        "temp_id": 541,
        "size": "381*-7268",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "202bcff812b872bdc3b35c1180cddedd",
        "bound_box": "1632,9544,2013,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1648,
                9544
            ],
            [
                2013,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google DeepMind",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 541,
        "temp_id": 542,
        "size": "365*-7268",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Google DeepMind[enabled,,]",
        "view_str": "f08490f4dc1456e50c91b5c8aa47c351",
        "bound_box": "1648,9544,2013,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google logo",
        "children": [
            544
        ],
        "focused": false,
        "bounds": [
            [
                2008,
                9544
            ],
            [
                2294,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 530,
        "temp_id": 543,
        "size": "286*-7268",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "031cde89017e9ebcc2b3e25bed6e95e4",
        "bound_box": "2008,9544,2294,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                2023,
                9544
            ],
            [
                2294,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google logo",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 543,
        "temp_id": 544,
        "size": "271*-7268",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Google logo[enabled,,]",
        "view_str": "f6649c2f91bcc2c941b2d0e23c880197",
        "bound_box": "2023,9544,2294,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            546
        ],
        "focused": false,
        "bounds": [
            [
                0,
                9681
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 103,
        "temp_id": 545,
        "size": "1084*-7405",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "67049e768ef110aa9225cda8bf46cb44",
        "bound_box": "0,9681,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            547
        ],
        "focused": false,
        "bounds": [
            [
                0,
                9681
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 545,
        "temp_id": 546,
        "size": "1084*-7405",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "103594fa3687b9eb010a0cb55c42e6a8",
        "bound_box": "0,9681,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 3,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            548,
            557,
            559
        ],
        "focused": false,
        "bounds": [
            [
                0,
                9681
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 546,
        "temp_id": 547,
        "size": "1084*-7405",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "af4a96a71350767ffda65ff752b99edf",
        "bound_box": "0,9681,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            549
        ],
        "focused": false,
        "bounds": [
            [
                0,
                9681
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 547,
        "temp_id": 548,
        "size": "1084*-7405",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "78957fc8d9d6bf28d42cd5753145ef6a",
        "bound_box": "0,9681,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            550,
            556
        ],
        "focused": false,
        "bounds": [
            [
                0,
                9681
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 548,
        "temp_id": 549,
        "size": "1084*-7405",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "9059e8fff283cdedad5a4073a983c285",
        "bound_box": "0,9681,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "About Google https://about.google › intl › ALL_us Browse All of Google's Products & Services",
        "children": [
            551,
            555
        ],
        "focused": false,
        "bounds": [
            [
                0,
                9681
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 549,
        "temp_id": 550,
        "size": "1084*-7405",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "9c5d4fd6cbc407fdd471ff6c769c1017",
        "bound_box": "0,9681,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            552
        ],
        "focused": false,
        "bounds": [
            [
                42,
                9720
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 550,
        "temp_id": 551,
        "size": "1000*-7444",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "14fc7afd7803359827765f00aca8214d",
        "bound_box": "42,9720,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            553,
            554
        ],
        "focused": false,
        "bounds": [
            [
                42,
                9720
            ],
            [
                937,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 551,
        "temp_id": 552,
        "size": "895*-7444",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "9826dd442ab9e59349c60ae7c517c893",
        "bound_box": "42,9720,937,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                147,
                9723
            ],
            [
                640,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "About Google",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 552,
        "temp_id": 553,
        "size": "493*-7447",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]About Google[enabled,,]",
        "view_str": "06acb0c5f002e7d282f527b5bf8c4382",
        "bound_box": "147,9723,640,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                147,
                9778
            ],
            [
                640,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "https://about.google › intl › ALL_us",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 552,
        "temp_id": 554,
        "size": "493*-7502",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]https://about.google › intl › ALL_us[enabled,,]",
        "view_str": "21c752d9405154cec132d7c107f70093",
        "bound_box": "147,9778,640,2276",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                9846
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Browse All of Google's Products & Services",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 550,
        "temp_id": 555,
        "size": "1000*-7570",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Browse All of Google's Products & Services[enabled,,]",
        "view_str": "b4fcc81d9e312d2359b21cf9530e44e7",
        "bound_box": "42,9846,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                952,
                9681
            ],
            [
                1081,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "About this result",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 549,
        "temp_id": 556,
        "size": "129*-7405",
        "signature": "[class]android.widget.Button[resource_id]None[visible]False[text]About this result[enabled,,]",
        "view_str": "1664121feb337e00ea038619161786d9",
        "bound_box": "952,9681,1081,2276",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            558
        ],
        "focused": false,
        "bounds": [
            [
                0,
                9998
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 547,
        "temp_id": 557,
        "size": "1084*-7722",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "63bf2cd5a03b0f0b3405663df6b2874f",
        "bound_box": "0,9998,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                10003
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Browse a list of Google products designed to help you work and play, stay organized, get answers, keep in touch, grow your business, and more.",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 557,
        "temp_id": 558,
        "size": "1000*-7727",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "878c281d0b3766ccf7fdaeef4dec05b1",
        "bound_box": "42,10003,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            560
        ],
        "focused": false,
        "bounds": [
            [
                0,
                10174
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 547,
        "temp_id": 559,
        "size": "1084*-7898",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "78957fc8d9d6bf28d42cd5753145ef6a",
        "bound_box": "0,10174,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            561
        ],
        "focused": false,
        "bounds": [
            [
                0,
                10192
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 559,
        "temp_id": 560,
        "size": "1084*-7916",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "115268acf822c3866e5eb7f133f34992",
        "bound_box": "0,10192,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            562
        ],
        "focused": false,
        "bounds": [
            [
                0,
                10192
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": true,
        "selected": false,
        "long_clickable": false,
        "parent": 560,
        "temp_id": 561,
        "size": "1084*-7916",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "571457d2e2dc2d5c0c79b5abc5f729af",
        "bound_box": "0,10192,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 7,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            563,
            565,
            567,
            569,
            571,
            573,
            575
        ],
        "focused": false,
        "bounds": [
            [
                0,
                10192
            ],
            [
                2483,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 561,
        "temp_id": 562,
        "size": "2483*-7916",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "fe2d825f68a3639c3f6b85583bce2e62",
        "bound_box": "0,10192,2483,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google Public Sector",
        "children": [
            564
        ],
        "focused": false,
        "bounds": [
            [
                42,
                10192
            ],
            [
                456,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 562,
        "temp_id": 563,
        "size": "414*-7916",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "7cc898d6d20eb354bacc5bc9afdc37a2",
        "bound_box": "42,10192,456,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                10192
            ],
            [
                456,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google Public Sector",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 563,
        "temp_id": 564,
        "size": "414*-7916",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Google Public Sector[enabled,,]",
        "view_str": "2df7be74408928c57f88d742a4537b62",
        "bound_box": "42,10192,456,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Commitments",
        "children": [
            566
        ],
        "focused": false,
        "bounds": [
            [
                451,
                10192
            ],
            [
                774,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 562,
        "temp_id": 565,
        "size": "323*-7916",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "ae64ddb68f33a7f4f4578175d626e7c3",
        "bound_box": "451,10192,774,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                469,
                10192
            ],
            [
                774,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Commitments",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 565,
        "temp_id": 566,
        "size": "305*-7916",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Commitments[enabled,,]",
        "view_str": "afbe78d49f2b9fb7029dbdcbc7de675c",
        "bound_box": "469,10192,774,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Stories",
        "children": [
            568
        ],
        "focused": false,
        "bounds": [
            [
                771,
                10192
            ],
            [
                973,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 562,
        "temp_id": 567,
        "size": "202*-7916",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "58f188e437cac16cf3ba915faf746a9e",
        "bound_box": "771,10192,973,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                784,
                10192
            ],
            [
                973,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Stories",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 567,
        "temp_id": 568,
        "size": "189*-7916",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Stories[enabled,,]",
        "view_str": "55fd62d4dcf00e804c2db301813bd8dd",
        "bound_box": "784,10192,973,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Designing Inclusive Products...",
        "children": [
            570
        ],
        "focused": false,
        "bounds": [
            [
                971,
                10192
            ],
            [
                1564,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 562,
        "temp_id": 569,
        "size": "593*-7916",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "1cf4e892197f6163d07b8a4e87b30a43",
        "bound_box": "971,10192,1564,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                987,
                10192
            ],
            [
                1564,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Designing Inclusive Products...",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 569,
        "temp_id": 570,
        "size": "577*-7916",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Designing Inclusive Products...[enabled,,]",
        "view_str": "24f71ef1a889c2875db21f11b23d28cf",
        "bound_box": "987,10192,1564,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Contact us",
        "children": [
            572
        ],
        "focused": false,
        "bounds": [
            [
                1561,
                10192
            ],
            [
                1827,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 562,
        "temp_id": 571,
        "size": "266*-7916",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "a4f8d86365910d7d471def6029d84c0e",
        "bound_box": "1561,10192,1827,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1577,
                10192
            ],
            [
                1827,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Contact us",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 571,
        "temp_id": 572,
        "size": "250*-7916",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Contact us[enabled,,]",
        "view_str": "94c98dfe5038583604ea9349d6417add",
        "bound_box": "1577,10192,1827,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Helpful products.",
        "children": [
            574
        ],
        "focused": false,
        "bounds": [
            [
                1821,
                10192
            ],
            [
                2194,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 562,
        "temp_id": 573,
        "size": "373*-7916",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "d2664f486add0bbbd6d33a1fb4b15efe",
        "bound_box": "1821,10192,2194,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1837,
                10192
            ],
            [
                2194,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Helpful products.",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 573,
        "temp_id": 574,
        "size": "357*-7916",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Helpful products.[enabled,,]",
        "view_str": "ad37c31ab644a37b0c8f0d336e109c5f",
        "bound_box": "1837,10192,2194,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Belonging",
        "children": [
            576
        ],
        "focused": false,
        "bounds": [
            [
                2189,
                10192
            ],
            [
                2441,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 562,
        "temp_id": 575,
        "size": "252*-7916",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "9b761763d4da5574f22b5814db3852ba",
        "bound_box": "2189,10192,2441,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                2205,
                10192
            ],
            [
                2441,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Belonging",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 575,
        "temp_id": 576,
        "size": "236*-7916",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Belonging[enabled,,]",
        "view_str": "8998ffd76237367ae1f8db968a79c35b",
        "bound_box": "2205,10192,2441,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                10326
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "bottomads",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 96,
        "temp_id": 577,
        "size": "1084*-8050",
        "signature": "[class]android.view.View[resource_id]bottomads[visible]False[text][enabled,,]",
        "view_str": "39a49333608466085f8ea30f38abe7ad",
        "bound_box": "0,10326,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]bottomads[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            579
        ],
        "focused": false,
        "bounds": [
            [
                0,
                10326
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "botstuff",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 96,
        "temp_id": 578,
        "size": "1084*-8050",
        "signature": "[class]android.view.View[resource_id]botstuff[visible]False[text][enabled,,]",
        "view_str": "acbf0e40f0d60e6cdf8696f198f1e004",
        "bound_box": "0,10326,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]botstuff[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 5,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            580,
            620,
            621,
            622,
            623
        ],
        "focused": false,
        "bounds": [
            [
                0,
                10326
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 578,
        "temp_id": 579,
        "size": "1084*-8050",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "c7071b6d68b45939fb98a49a7bcb9ba7",
        "bound_box": "0,10326,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            581
        ],
        "focused": false,
        "bounds": [
            [
                0,
                10326
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "bres",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 579,
        "temp_id": 580,
        "size": "1084*-8050",
        "signature": "[class]android.view.View[resource_id]bres[visible]False[text][enabled,,]",
        "view_str": "5955323f74da174972a37356c33dc40a",
        "bound_box": "0,10326,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]bres[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 12,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            582,
            585,
            590,
            591,
            596,
            597,
            602,
            603,
            608,
            609,
            614,
            615
        ],
        "focused": false,
        "bounds": [
            [
                0,
                10326
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 580,
        "temp_id": 581,
        "size": "1084*-8050",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "ba407c4ca55ed0afa35042f0366bb8e4",
        "bound_box": "0,10326,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            583,
            584
        ],
        "focused": false,
        "bounds": [
            [
                0,
                10326
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 581,
        "temp_id": 582,
        "size": "1084*-8050",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "eef4237f8c2afb76bcbba41ba4767c13",
        "bound_box": "0,10326,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                10368
            ],
            [
                1010,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "People also search for",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 582,
        "temp_id": 583,
        "size": "968*-8092",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]People also search for[enabled,,]",
        "view_str": "f565aed954dcd7629cf072cecf069dc9",
        "bound_box": "42,10368,1010,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                952,
                10326
            ],
            [
                1081,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "About this result",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 582,
        "temp_id": 584,
        "size": "129*-8050",
        "signature": "[class]android.widget.Button[resource_id]None[visible]False[text]About this result[enabled,,]",
        "view_str": "8c679f1fe7aa991c503c09d2523b756b",
        "bound_box": "952,10326,1081,2276",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            586
        ],
        "focused": false,
        "bounds": [
            [
                42,
                10479
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": "2-0yZ-jtAcyGptQPofi-iA8__156",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 581,
        "temp_id": 585,
        "size": "1000*-8203",
        "signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__156[visible]False[text][enabled,,]",
        "view_str": "4a54524a42bef3e3dce50b082150d705",
        "bound_box": "42,10479,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__156[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            587
        ],
        "focused": false,
        "bounds": [
            [
                42,
                10479
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 585,
        "temp_id": 586,
        "size": "1000*-8203",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "83f6b77ca3dc9e80a02a23a52cf24675",
        "bound_box": "42,10479,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google Play",
        "children": [
            588,
            589
        ],
        "focused": false,
        "bounds": [
            [
                42,
                10479
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 586,
        "temp_id": 587,
        "size": "1000*-8203",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "9c30c2425cd8df63fb917bfe93c810f9",
        "bound_box": "42,10479,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                10531
            ],
            [
                916,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google Play",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 587,
        "temp_id": 588,
        "size": "874*-8255",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Google Play[enabled,,]",
        "view_str": "426f8b67076c780c261d9990ef96b649",
        "bound_box": "42,10531,916,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                968,
                10531
            ],
            [
                1023,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.widget.Image",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 587,
        "temp_id": 589,
        "size": "55*-8255",
        "signature": "[class]android.widget.Image[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "6a7e7bbbe8364f68527b01398984a69a",
        "bound_box": "968,10531,1023,2276",
        "content_free_signature": "[class]android.widget.Image[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                10636
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 581,
        "temp_id": 590,
        "size": "1000*-8360",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "2c789f651be2edaf384fe1519307e772",
        "bound_box": "42,10636,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            592
        ],
        "focused": false,
        "bounds": [
            [
                42,
                10639
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": "2-0yZ-jtAcyGptQPofi-iA8__157",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 581,
        "temp_id": 591,
        "size": "1000*-8363",
        "signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__157[visible]False[text][enabled,,]",
        "view_str": "5b310051284d82fa6614c418158c27f5",
        "bound_box": "42,10639,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__157[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            593
        ],
        "focused": false,
        "bounds": [
            [
                42,
                10639
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 591,
        "temp_id": 592,
        "size": "1000*-8363",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "db2cf12a0fae2d071c214b679802b6a8",
        "bound_box": "42,10639,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google sign in",
        "children": [
            594,
            595
        ],
        "focused": false,
        "bounds": [
            [
                42,
                10639
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 592,
        "temp_id": 593,
        "size": "1000*-8363",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "d0a8398de3c45329fa26f6cba2001861",
        "bound_box": "42,10639,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                10691
            ],
            [
                916,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google sign in",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 593,
        "temp_id": 594,
        "size": "874*-8415",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Google sign in[enabled,,]",
        "view_str": "91ec26af735733a27dd86d4c67fdb19a",
        "bound_box": "42,10691,916,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                968,
                10691
            ],
            [
                1023,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.widget.Image",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 593,
        "temp_id": 595,
        "size": "55*-8415",
        "signature": "[class]android.widget.Image[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "0f002b7497beb28d7f2d2f701134a608",
        "bound_box": "968,10691,1023,2276",
        "content_free_signature": "[class]android.widget.Image[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                10796
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 581,
        "temp_id": 596,
        "size": "1000*-8520",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "2c789f651be2edaf384fe1519307e772",
        "bound_box": "42,10796,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            598
        ],
        "focused": false,
        "bounds": [
            [
                42,
                10799
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": "2-0yZ-jtAcyGptQPofi-iA8__158",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 581,
        "temp_id": 597,
        "size": "1000*-8523",
        "signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__158[visible]False[text][enabled,,]",
        "view_str": "f6381080e0c6d183e2b12ca5796a852d",
        "bound_box": "42,10799,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__158[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            599
        ],
        "focused": false,
        "bounds": [
            [
                42,
                10799
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 597,
        "temp_id": 598,
        "size": "1000*-8523",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "57061f479928cbb6eabc455778b6a671",
        "bound_box": "42,10799,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google Chrome",
        "children": [
            600,
            601
        ],
        "focused": false,
        "bounds": [
            [
                42,
                10799
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 598,
        "temp_id": 599,
        "size": "1000*-8523",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "734f0b49fe9e4b4bae0a04629a5ec341",
        "bound_box": "42,10799,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                10851
            ],
            [
                916,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google Chrome",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 599,
        "temp_id": 600,
        "size": "874*-8575",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Google Chrome[enabled,,]",
        "view_str": "2bc4b7627f74be689669fd0869876534",
        "bound_box": "42,10851,916,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                968,
                10851
            ],
            [
                1023,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.widget.Image",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 599,
        "temp_id": 601,
        "size": "55*-8575",
        "signature": "[class]android.widget.Image[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "b81397200a3898c7faebbaf75e0c5be8",
        "bound_box": "968,10851,1023,2276",
        "content_free_signature": "[class]android.widget.Image[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                10956
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 581,
        "temp_id": 602,
        "size": "1000*-8680",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "2c789f651be2edaf384fe1519307e772",
        "bound_box": "42,10956,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            604
        ],
        "focused": false,
        "bounds": [
            [
                42,
                10959
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": "2-0yZ-jtAcyGptQPofi-iA8__159",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 581,
        "temp_id": 603,
        "size": "1000*-8683",
        "signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__159[visible]False[text][enabled,,]",
        "view_str": "f6734963e51c13e451f066d9b844dd5c",
        "bound_box": "42,10959,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__159[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            605
        ],
        "focused": false,
        "bounds": [
            [
                42,
                10959
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 603,
        "temp_id": 604,
        "size": "1000*-8683",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "c28329d9f045ea80c98f65ac1fd50bbd",
        "bound_box": "42,10959,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google Pay",
        "children": [
            606,
            607
        ],
        "focused": false,
        "bounds": [
            [
                42,
                10959
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 604,
        "temp_id": 605,
        "size": "1000*-8683",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "bd93ef2ef71b7f5f3f86adbd39f89ce7",
        "bound_box": "42,10959,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                11011
            ],
            [
                916,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google Pay",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 605,
        "temp_id": 606,
        "size": "874*-8735",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Google Pay[enabled,,]",
        "view_str": "0448cd2592b33e42210b2f2821c6a821",
        "bound_box": "42,11011,916,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                968,
                11011
            ],
            [
                1023,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.widget.Image",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 605,
        "temp_id": 607,
        "size": "55*-8735",
        "signature": "[class]android.widget.Image[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "46adcd1095375aa07ebcd692f5b592da",
        "bound_box": "968,11011,1023,2276",
        "content_free_signature": "[class]android.widget.Image[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                11116
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 581,
        "temp_id": 608,
        "size": "1000*-8840",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "2c789f651be2edaf384fe1519307e772",
        "bound_box": "42,11116,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            610
        ],
        "focused": false,
        "bounds": [
            [
                42,
                11119
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": "2-0yZ-jtAcyGptQPofi-iA8__160",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 581,
        "temp_id": 609,
        "size": "1000*-8843",
        "signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__160[visible]False[text][enabled,,]",
        "view_str": "5feb14da44f056fa604aa185943ae723",
        "bound_box": "42,11119,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__160[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            611
        ],
        "focused": false,
        "bounds": [
            [
                42,
                11119
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 609,
        "temp_id": 610,
        "size": "1000*-8843",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "667a6211ef4b25f6ba7b9395b4074025",
        "bound_box": "42,11119,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google history",
        "children": [
            612,
            613
        ],
        "focused": false,
        "bounds": [
            [
                42,
                11119
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 610,
        "temp_id": 611,
        "size": "1000*-8843",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "80356b38973dcb60fab68db795ccb352",
        "bound_box": "42,11119,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                11172
            ],
            [
                916,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google history",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 611,
        "temp_id": 612,
        "size": "874*-8896",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Google history[enabled,,]",
        "view_str": "3c2de90357f2f6cc179d870e956bdc7c",
        "bound_box": "42,11172,916,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                968,
                11172
            ],
            [
                1023,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.widget.Image",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 611,
        "temp_id": 613,
        "size": "55*-8896",
        "signature": "[class]android.widget.Image[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "821ab69e2441f2f1d566a6e00cb0d4fb",
        "bound_box": "968,11172,1023,2276",
        "content_free_signature": "[class]android.widget.Image[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                11277
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 581,
        "temp_id": 614,
        "size": "1000*-9001",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "2c789f651be2edaf384fe1519307e772",
        "bound_box": "42,11277,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            616
        ],
        "focused": false,
        "bounds": [
            [
                42,
                11279
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": "2-0yZ-jtAcyGptQPofi-iA8__161",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 581,
        "temp_id": 615,
        "size": "1000*-9003",
        "signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__161[visible]False[text][enabled,,]",
        "view_str": "510f5c85819a8d8c17300feb922ed51e",
        "bound_box": "42,11279,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]2-0yZ-jtAcyGptQPofi-iA8__161[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            617
        ],
        "focused": false,
        "bounds": [
            [
                42,
                11279
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 615,
        "temp_id": 616,
        "size": "1000*-9003",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "8ec913d48c76751716caa3761f98e88a",
        "bound_box": "42,11279,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Google Play Store",
        "children": [
            618,
            619
        ],
        "focused": false,
        "bounds": [
            [
                42,
                11279
            ],
            [
                1042,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 616,
        "temp_id": 617,
        "size": "1000*-9003",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "04b8297d235a0b1960421cd284df3ce9",
        "bound_box": "42,11279,1042,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                42,
                11332
            ],
            [
                916,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Google Play Store",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 617,
        "temp_id": 618,
        "size": "874*-9056",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Google Play Store[enabled,,]",
        "view_str": "2ba03ddde1e0c2f5b9f71ded5cdde272",
        "bound_box": "42,11332,916,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                968,
                11332
            ],
            [
                1023,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.widget.Image",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 617,
        "temp_id": 619,
        "size": "55*-9056",
        "signature": "[class]android.widget.Image[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "312c3e02e65acd1e3f82878c3fc8a654",
        "bound_box": "968,11332,1023,2276",
        "content_free_signature": "[class]android.widget.Image[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                11463
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "arc-srp_2-0yZ-jtAcyGptQPofi-iA8_1",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 579,
        "temp_id": 620,
        "size": "1084*-9187",
        "signature": "[class]android.view.View[resource_id]arc-srp_2-0yZ-jtAcyGptQPofi-iA8_1[visible]False[text][enabled,,]",
        "view_str": "d52d724953e40ed902a31f4310d6ff80",
        "bound_box": "0,11463,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]arc-srp_2-0yZ-jtAcyGptQPofi-iA8_1[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                11515
            ],
            [
                5,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Page Navigation",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 579,
        "temp_id": 621,
        "size": "5*-9239",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Page Navigation[enabled,,]",
        "view_str": "2ffd1cb011d0b00be3ab3ffa34a9e923",
        "bound_box": "0,11515,5,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                11515
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "More search results",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 579,
        "temp_id": 622,
        "size": "1084*-9239",
        "signature": "[class]android.widget.Button[resource_id]None[visible]False[text]More search results[enabled,,]",
        "view_str": "87086434428b53167fb7a479b20cad36",
        "bound_box": "0,11515,1084,2276",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            624
        ],
        "focused": false,
        "bounds": [
            [
                0,
                11959
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 579,
        "temp_id": 623,
        "size": "1084*-9683",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "ebf09012cc22a58d47fc2c49edb8c615",
        "bound_box": "0,11959,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                11673
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 623,
        "temp_id": 624,
        "size": "1084*-9397",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "d0ff2e737614e9cb59ef46f9399f1ccf",
        "bound_box": "0,11673,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                11683
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 96,
        "temp_id": 625,
        "size": "1084*-9407",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "6f38360104f946ec9e396e9a5f157084",
        "bound_box": "0,11683,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                2275
            ],
            [
                1084,
                2275
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 33,
        "temp_id": 626,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "1d64df32b47d1ad640421a476c1e93c2",
        "bound_box": "0,2275,1084,2275",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            628
        ],
        "focused": false,
        "bounds": [
            [
                0,
                2275
            ],
            [
                1084,
                2275
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 33,
        "temp_id": 627,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "c1bb2932cc410a20a8b50d66f5e7d2e0",
        "bound_box": "0,2275,1084,2275",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                2275
            ],
            [
                1084,
                2275
            ]
        ],
        "resource_id": "rNi7Zc",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 627,
        "temp_id": 628,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]rNi7Zc[visible]False[text][enabled,,]",
        "view_str": "57e3150a123550d5c470cc4c77912d4e",
        "bound_box": "0,2275,1084,2275",
        "content_free_signature": "[class]android.view.View[resource_id]rNi7Zc[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            630
        ],
        "focused": false,
        "bounds": [
            [
                0,
                2275
            ],
            [
                1084,
                2275
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 33,
        "temp_id": 629,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "c1bb2932cc410a20a8b50d66f5e7d2e0",
        "bound_box": "0,2275,1084,2275",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                2275
            ],
            [
                1084,
                2275
            ]
        ],
        "resource_id": "rNi7Zc",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 629,
        "temp_id": 630,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]rNi7Zc[visible]False[text][enabled,,]",
        "view_str": "57e3150a123550d5c470cc4c77912d4e",
        "bound_box": "0,2275,1084,2275",
        "content_free_signature": "[class]android.view.View[resource_id]rNi7Zc[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            632
        ],
        "focused": false,
        "bounds": [
            [
                0,
                2275
            ],
            [
                1084,
                2275
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 33,
        "temp_id": 631,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "c1bb2932cc410a20a8b50d66f5e7d2e0",
        "bound_box": "0,2275,1084,2275",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                2275
            ],
            [
                1084,
                2275
            ]
        ],
        "resource_id": "rNi7Zc",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 631,
        "temp_id": 632,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]rNi7Zc[visible]False[text][enabled,,]",
        "view_str": "57e3150a123550d5c470cc4c77912d4e",
        "bound_box": "0,2275,1084,2275",
        "content_free_signature": "[class]android.view.View[resource_id]rNi7Zc[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            634
        ],
        "focused": false,
        "bounds": [
            [
                0,
                2275
            ],
            [
                1084,
                2275
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 33,
        "temp_id": 633,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "c1bb2932cc410a20a8b50d66f5e7d2e0",
        "bound_box": "0,2275,1084,2275",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                2275
            ],
            [
                1084,
                2275
            ]
        ],
        "resource_id": "rNi7Zc",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 633,
        "temp_id": 634,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]rNi7Zc[visible]False[text][enabled,,]",
        "view_str": "57e3150a123550d5c470cc4c77912d4e",
        "bound_box": "0,2275,1084,2275",
        "content_free_signature": "[class]android.view.View[resource_id]rNi7Zc[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            636
        ],
        "focused": false,
        "bounds": [
            [
                0,
                11683
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "sfooter",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 33,
        "temp_id": 635,
        "size": "1084*-9407",
        "signature": "[class]android.view.View[resource_id]sfooter[visible]False[text][enabled,,]",
        "view_str": "686b59dbb59d01753541ed5f376c8fac",
        "bound_box": "0,11683,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]sfooter[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            637,
            638
        ],
        "focused": false,
        "bounds": [
            [
                0,
                11683
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "bfb_2-0yZ-jtAcyGptQPofi-iA8_1",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 635,
        "temp_id": 636,
        "size": "1084*-9407",
        "signature": "[class]android.view.View[resource_id]bfb_2-0yZ-jtAcyGptQPofi-iA8_1[visible]False[text][enabled,,]",
        "view_str": "baf64c63ec363924c0ddb1a9493242c6",
        "bound_box": "0,11683,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]bfb_2-0yZ-jtAcyGptQPofi-iA8_1[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                11683
            ],
            [
                5,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Footer Links",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 636,
        "temp_id": 637,
        "size": "5*-9407",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]Footer Links[enabled,,]",
        "view_str": "e579ed91c757f260a5cb3123325ca7bc",
        "bound_box": "0,11683,5,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 3,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            639,
            646,
            653
        ],
        "focused": false,
        "bounds": [
            [
                0,
                11683
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "fbar",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 636,
        "temp_id": 638,
        "size": "1084*-9407",
        "signature": "[class]android.view.View[resource_id]fbar[visible]False[text][enabled,,]",
        "view_str": "ab67ba7a073f2419158b5324e2318b3f",
        "bound_box": "0,11683,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]fbar[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 3,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            640,
            641,
            644
        ],
        "focused": false,
        "bounds": [
            [
                0,
                11725
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "swml",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 638,
        "temp_id": 639,
        "size": "1084*-9449",
        "signature": "[class]android.view.View[resource_id]swml[visible]False[text][enabled,,]",
        "view_str": "eca33570da6cc6990aa35a915b4fbecd",
        "bound_box": "0,11725,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]swml[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                147,
                11757
            ],
            [
                934,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "94043, Mountain View, CA - From your device",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 639,
        "temp_id": 640,
        "size": "787*-9481",
        "signature": "[class]android.widget.Button[resource_id]None[visible]False[text]94043, Mountain View, CA - From your device[enabled,,]",
        "view_str": "96b4ec946dfc7cd134d37769ef5e34e8",
        "bound_box": "147,11757,934,2276",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            642
        ],
        "focused": false,
        "bounds": [
            [
                147,
                12096
            ],
            [
                934,
                2276
            ]
        ],
        "resource_id": "tsuid_2-0yZ-jtAcyGptQPofi-iA8_12",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 639,
        "temp_id": 641,
        "size": "787*-9820",
        "signature": "[class]android.view.View[resource_id]tsuid_2-0yZ-jtAcyGptQPofi-iA8_12[visible]False[text][enabled,,]",
        "view_str": "3490f0135d60a357e36e2fcc6ba8f4f9",
        "bound_box": "147,12096,934,2276",
        "content_free_signature": "[class]android.view.View[resource_id]tsuid_2-0yZ-jtAcyGptQPofi-iA8_12[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            643
        ],
        "focused": false,
        "bounds": [
            [
                147,
                12096
            ],
            [
                934,
                2276
            ]
        ],
        "resource_id": "ow22",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 641,
        "temp_id": 642,
        "size": "787*-9820",
        "signature": "[class]android.view.View[resource_id]ow22[visible]False[text][enabled,,]",
        "view_str": "8fe1f89417ec260152c9d99c8ebc0b09",
        "bound_box": "147,12096,934,2276",
        "content_free_signature": "[class]android.view.View[resource_id]ow22[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                210
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_16",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 642,
        "temp_id": 643,
        "size": "1084*2066",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_16[visible]True[text][enabled,,]",
        "view_str": "52a4f79ad1935baeea4eda3fa5301d8c",
        "bound_box": "0,210,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_16[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            645
        ],
        "focused": false,
        "bounds": [
            [
                0,
                11830
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 639,
        "temp_id": 644,
        "size": "1084*-9554",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "2d4fdc70c4115c2e11b6399d23fe23cd",
        "bound_box": "0,11830,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                409,
                11854
            ],
            [
                672,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Update location",
        "class": "android.widget.Button",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 644,
        "temp_id": 645,
        "size": "263*-9578",
        "signature": "[class]android.widget.Button[resource_id]None[visible]False[text]Update location[enabled,,]",
        "view_str": "395cbf4edd6ddd6b6645e9703188dc66",
        "bound_box": "409,11854,672,2276",
        "content_free_signature": "[class]android.widget.Button[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 3,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            647,
            649,
            651
        ],
        "focused": false,
        "bounds": [
            [
                -73,
                11935
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 638,
        "temp_id": 646,
        "size": "1157*-9659",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "05269ea2156ad574dfbe12c9b84c8939",
        "bound_box": "-73,11935,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Dark theme: off",
        "children": [
            648
        ],
        "focused": false,
        "bounds": [
            [
                154,
                11935
            ],
            [
                480,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 646,
        "temp_id": 647,
        "size": "326*-9659",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "2be5911a40897132d980328dd250a1b7",
        "bound_box": "154,11935,480,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                225,
                11959
            ],
            [
                480,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Dark theme: off",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 647,
        "temp_id": 648,
        "size": "255*-9683",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]Dark theme: off[enabled,,]",
        "view_str": "bca7173eb4ba9e2f0004cf8153dd2a15",
        "bound_box": "225,11959,480,2276",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Help",
        "children": [
            650
        ],
        "focused": false,
        "bounds": [
            [
                477,
                11935
            ],
            [
                627,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 646,
        "temp_id": 649,
        "size": "150*-9659",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "06ee0a3d0eb8d436dd95f1564d720da2",
        "bound_box": "477,11935,627,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                548,
                11959
            ],
            [
                627,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Help",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 649,
        "temp_id": 650,
        "size": "79*-9683",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]Help[enabled,,]",
        "view_str": "90b161c77a8a7ad52fbfb39eb7d3a21e",
        "bound_box": "548,11959,627,2276",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Feedback",
        "children": [
            652
        ],
        "focused": false,
        "bounds": [
            [
                624,
                11935
            ],
            [
                855,
                2276
            ]
        ],
        "resource_id": "dk2qOd",
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 646,
        "temp_id": 651,
        "size": "231*-9659",
        "signature": "[class]android.view.View[resource_id]dk2qOd[visible]False[text]None[enabled,,]",
        "view_str": "9905dab775651de49d00d53ee307d378",
        "bound_box": "624,11935,855,2276",
        "content_free_signature": "[class]android.view.View[resource_id]dk2qOd[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                695,
                11959
            ],
            [
                855,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Feedback",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 651,
        "temp_id": 652,
        "size": "160*-9683",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]Feedback[enabled,,]",
        "view_str": "d504f25e70276612c1951bccc9e8693f",
        "bound_box": "695,11959,855,2276",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            654,
            656
        ],
        "focused": false,
        "bounds": [
            [
                -73,
                12027
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 638,
        "temp_id": 653,
        "size": "1157*-9751",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "b72c077b72b9b0445b628ea371fb683d",
        "bound_box": "-73,12027,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Privacy",
        "children": [
            655
        ],
        "focused": false,
        "bounds": [
            [
                322,
                12027
            ],
            [
                514,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 653,
        "temp_id": 654,
        "size": "192*-9751",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "6cffc8fcbae0dfdc17d64ac63fed3072",
        "bound_box": "322,12027,514,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                393,
                12051
            ],
            [
                514,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Privacy",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 654,
        "temp_id": 655,
        "size": "121*-9775",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]Privacy[enabled,,]",
        "view_str": "9d521ee32df3c186fa2c4b0c4d3b9350",
        "bound_box": "393,12051,514,2276",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Terms",
        "children": [
            657
        ],
        "focused": false,
        "bounds": [
            [
                511,
                12027
            ],
            [
                690,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 653,
        "temp_id": 656,
        "size": "179*-9751",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "a5801fbe672bb61d9b46ccc4464b6571",
        "bound_box": "511,12027,690,2276",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                582,
                12051
            ],
            [
                690,
                2276
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "Terms",
        "class": "android.widget.TextView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 656,
        "temp_id": 657,
        "size": "108*-9775",
        "signature": "[class]android.widget.TextView[resource_id]None[visible]False[text]Terms[enabled,,]",
        "view_str": "f43433ad719243aa8ba9c7b94d3b64a3",
        "bound_box": "582,12051,690,2276",
        "content_free_signature": "[class]android.widget.TextView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            659
        ],
        "focused": false,
        "bounds": [
            [
                0,
                12190
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_36",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 32,
        "temp_id": 658,
        "size": "1084*-9914",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_36[visible]False[text][enabled,,]",
        "view_str": "6b63d7ee89dfade55857f51308e37cfb",
        "bound_box": "0,12190,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_36[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                12190
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "_2-0yZ-jtAcyGptQPofi-iA8_39",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 658,
        "temp_id": 659,
        "size": "1084*-9914",
        "signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_39[visible]False[text][enabled,,]",
        "view_str": "8633f81f79f1588ea03e292c56f479fc",
        "bound_box": "0,12190,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]_2-0yZ-jtAcyGptQPofi-iA8_39[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            661
        ],
        "focused": false,
        "bounds": [
            [
                0,
                12190
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "TWfxFb",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 11,
        "temp_id": 660,
        "size": "1084*-9914",
        "signature": "[class]android.view.View[resource_id]TWfxFb[visible]False[text][enabled,,]",
        "view_str": "046c255fd472d25fc4ce405460bc6125",
        "bound_box": "0,12190,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]TWfxFb[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                12190
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "QPwIld",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 660,
        "temp_id": 661,
        "size": "1084*-9914",
        "signature": "[class]android.view.View[resource_id]QPwIld[visible]False[text][enabled,,]",
        "view_str": "8088a6382e205d445dd118b6e67a644c",
        "bound_box": "0,12190,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]QPwIld[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                12190
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "gws-plugins-collections-tray__save-components-async",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 11,
        "temp_id": 662,
        "size": "1084*-9914",
        "signature": "[class]android.view.View[resource_id]gws-plugins-collections-tray__save-components-async[visible]False[text][enabled,,]",
        "view_str": "7c3334b7e832d1b674b9e11d67676cd8",
        "bound_box": "0,12190,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]gws-plugins-collections-tray__save-components-async[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            664
        ],
        "focused": false,
        "bounds": [
            [
                0,
                12190
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "lfootercc",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 11,
        "temp_id": 663,
        "size": "1084*-9914",
        "signature": "[class]android.view.View[resource_id]lfootercc[visible]False[text][enabled,,]",
        "view_str": "ddcd66a4a44a14db1dd53b0750ce521f",
        "bound_box": "0,12190,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]lfootercc[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                12190
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "dbg_",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 663,
        "temp_id": 664,
        "size": "1084*-9914",
        "signature": "[class]android.view.View[resource_id]dbg_[visible]False[text][enabled,,]",
        "view_str": "2cd82fc713793648cd197b512bd2403f",
        "bound_box": "0,12190,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]dbg_[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                210
            ],
            [
                1084,
                2276
            ]
        ],
        "resource_id": "sZmt3b",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 11,
        "temp_id": 665,
        "size": "1084*2066",
        "signature": "[class]android.view.View[resource_id]sZmt3b[visible]True[text][enabled,,]",
        "view_str": "7eb4b68ff126234a7d1e963859181c7c",
        "bound_box": "0,210,1084,2276",
        "content_free_signature": "[class]android.view.View[resource_id]sZmt3b[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 7,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            667,
            668,
            669,
            670,
            671,
            672,
            673
        ],
        "focused": false,
        "bounds": [
            [
                0,
                2275
            ],
            [
                1084,
                2275
            ]
        ],
        "resource_id": "snbc",
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 11,
        "temp_id": 666,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]snbc[visible]False[text][enabled,,]",
        "view_str": "a5f10c1cf015ae1c361535dc7e8a5a9b",
        "bound_box": "0,2275,1084,2275",
        "content_free_signature": "[class]android.view.View[resource_id]snbc[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                2275
            ],
            [
                1084,
                2275
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 666,
        "temp_id": 667,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "0b3e80e76ca1e194b8a4ed2e6c9546b4",
        "bound_box": "0,2275,1084,2275",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                2275
            ],
            [
                1084,
                2275
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 666,
        "temp_id": 668,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "0b3e80e76ca1e194b8a4ed2e6c9546b4",
        "bound_box": "0,2275,1084,2275",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                2275
            ],
            [
                1084,
                2275
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 666,
        "temp_id": 669,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "0b3e80e76ca1e194b8a4ed2e6c9546b4",
        "bound_box": "0,2275,1084,2275",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                2275
            ],
            [
                1084,
                2275
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 666,
        "temp_id": 670,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "0b3e80e76ca1e194b8a4ed2e6c9546b4",
        "bound_box": "0,2275,1084,2275",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                2275
            ],
            [
                1084,
                2275
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 666,
        "temp_id": 671,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "0b3e80e76ca1e194b8a4ed2e6c9546b4",
        "bound_box": "0,2275,1084,2275",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                2275
            ],
            [
                1084,
                2275
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 666,
        "temp_id": 672,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "0b3e80e76ca1e194b8a4ed2e6c9546b4",
        "bound_box": "0,2275,1084,2275",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                2275
            ],
            [
                1084,
                2275
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": "",
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 666,
        "temp_id": 673,
        "size": "1084*0",
        "signature": "[class]android.view.View[resource_id]None[visible]False[text][enabled,,]",
        "view_str": "0b3e80e76ca1e194b8a4ed2e6c9546b4",
        "bound_box": "0,2275,1084,2275",
        "content_free_signature": "[class]android.view.View[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            675
        ],
        "focused": false,
        "bounds": [
            [
                0,
                63
            ],
            [
                1080,
                231
            ]
        ],
        "resource_id": "com.android.chrome:id/control_container",
        "checked": false,
        "text": null,
        "class": "android.widget.FrameLayout",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 5,
        "temp_id": 674,
        "size": "1080*168",
        "signature": "[class]android.widget.FrameLayout[resource_id]com.android.chrome:id/control_container[visible]True[text]None[enabled,,]",
        "view_str": "84f2d970ffe1f230d949ea02c73e9ae6",
        "bound_box": "0,63,1080,231",
        "content_free_signature": "[class]android.widget.FrameLayout[resource_id]com.android.chrome:id/control_container[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            676,
            687
        ],
        "focused": false,
        "bounds": [
            [
                0,
                63
            ],
            [
                1080,
                231
            ]
        ],
        "resource_id": "com.android.chrome:id/toolbar_container",
        "checked": false,
        "text": null,
        "class": "android.widget.FrameLayout",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 674,
        "temp_id": 675,
        "size": "1080*168",
        "signature": "[class]android.widget.FrameLayout[resource_id]com.android.chrome:id/toolbar_container[visible]True[text]None[enabled,,]",
        "view_str": "c825723a7abc20956466ebc56aca1215",
        "bound_box": "0,63,1080,231",
        "content_free_signature": "[class]android.widget.FrameLayout[resource_id]com.android.chrome:id/toolbar_container[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 3,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            677,
            678,
            682
        ],
        "focused": false,
        "bounds": [
            [
                0,
                63
            ],
            [
                1080,
                210
            ]
        ],
        "resource_id": "com.android.chrome:id/toolbar",
        "checked": false,
        "text": null,
        "class": "android.widget.FrameLayout",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 675,
        "temp_id": 676,
        "size": "1080*147",
        "signature": "[class]android.widget.FrameLayout[resource_id]com.android.chrome:id/toolbar[visible]True[text]None[enabled,,]",
        "view_str": "45b12259e7783e16553a8be75d893458",
        "bound_box": "0,63,1080,210",
        "content_free_signature": "[class]android.widget.FrameLayout[resource_id]com.android.chrome:id/toolbar[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Home",
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                63
            ],
            [
                126,
                210
            ]
        ],
        "resource_id": "com.android.chrome:id/home_button",
        "checked": false,
        "text": null,
        "class": "android.widget.ImageButton",
        "scrollable": false,
        "selected": false,
        "long_clickable": true,
        "parent": 676,
        "temp_id": 677,
        "size": "126*147",
        "signature": "[class]android.widget.ImageButton[resource_id]com.android.chrome:id/home_button[visible]True[text]None[enabled,,]",
        "view_str": "fd62abe918f585b3b0c24e9410aa2990",
        "bound_box": "0,63,126,210",
        "content_free_signature": "[class]android.widget.ImageButton[resource_id]com.android.chrome:id/home_button[visible]True",
        "allowed_actions": [
            "touch",
            "long_touch"
        ],
        "status": [],
        "local_id": "82",
        "full_desc": "<button alt='Home' bound_box=0,63,126,210></button>",
        "desc": "<button alt='Home' bound_box=0,63,126,210></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            679,
            681
        ],
        "focused": false,
        "bounds": [
            [
                126,
                63
            ],
            [
                828,
                210
            ]
        ],
        "resource_id": "com.android.chrome:id/location_bar",
        "checked": false,
        "text": null,
        "class": "android.widget.FrameLayout",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 676,
        "temp_id": 678,
        "size": "702*147",
        "signature": "[class]android.widget.FrameLayout[resource_id]com.android.chrome:id/location_bar[visible]True[text]None[enabled,,]",
        "view_str": "89e84e55b93e03b8db2f8feec2813800",
        "bound_box": "126,63,828,210",
        "content_free_signature": "[class]android.widget.FrameLayout[resource_id]com.android.chrome:id/location_bar[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            680
        ],
        "focused": false,
        "bounds": [
            [
                147,
                63
            ],
            [
                220,
                210
            ]
        ],
        "resource_id": "com.android.chrome:id/location_bar_status",
        "checked": false,
        "text": null,
        "class": "android.widget.LinearLayout",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 678,
        "temp_id": 679,
        "size": "73*147",
        "signature": "[class]android.widget.LinearLayout[resource_id]com.android.chrome:id/location_bar_status[visible]True[text]None[enabled,,]",
        "view_str": "ff05eabb5b32eb775f9cdea1efc4bfbb",
        "bound_box": "147,63,220,210",
        "content_free_signature": "[class]android.widget.LinearLayout[resource_id]com.android.chrome:id/location_bar_status[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Connection is secure. Site information",
        "children": [],
        "focused": false,
        "bounds": [
            [
                147,
                63
            ],
            [
                210,
                210
            ]
        ],
        "resource_id": "com.android.chrome:id/location_bar_status_icon",
        "checked": false,
        "text": null,
        "class": "android.widget.ImageButton",
        "scrollable": false,
        "selected": false,
        "long_clickable": true,
        "parent": 679,
        "temp_id": 680,
        "size": "63*147",
        "signature": "[class]android.widget.ImageButton[resource_id]com.android.chrome:id/location_bar_status_icon[visible]True[text]None[enabled,,]",
        "view_str": "30e3fde07599e5e2c7e14f77de5616f2",
        "bound_box": "147,63,210,210",
        "content_free_signature": "[class]android.widget.ImageButton[resource_id]com.android.chrome:id/location_bar_status_icon[visible]True",
        "allowed_actions": [
            "touch",
            "long_touch"
        ],
        "status": [],
        "local_id": "83",
        "full_desc": "<button alt='Connection is secure. Site information' bound_box=147,63,210,210></button>",
        "desc": "<button alt='Connection is secure. Site information' bound_box=147,63,210,210></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": true,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                220,
                71
            ],
            [
                807,
                202
            ]
        ],
        "resource_id": "com.android.chrome:id/url_bar",
        "checked": false,
        "text": "google.com.hk/search?gs_ssp=eJzj4tTP1TcwMU02T1JgNGB0YPBiS8_PT89JBQBASQXT&q=google&oq&aqs=chrome.3.69i58j35i39i362i523l2j46i39i199i362i465i523j35i39i362i523l3...6.-1j0j4&client=ms-unknown&sourceid=chrome-mobile&ie=UTF-8&gfe_rd=mr&pli=1",
        "class": "android.widget.EditText",
        "scrollable": false,
        "selected": false,
        "long_clickable": true,
        "parent": 678,
        "temp_id": 681,
        "size": "587*131",
        "signature": "[class]android.widget.EditText[resource_id]com.android.chrome:id/url_bar[visible]True[text]None[enabled,,]",
        "view_str": "ecc133c7d67accd8fd991ae9d6da3cf3",
        "bound_box": "220,71,807,202",
        "content_free_signature": "[class]android.widget.EditText[resource_id]com.android.chrome:id/url_bar[visible]True",
        "allowed_actions": [
            "touch",
            "set_text",
            "long_touch"
        ],
        "status": [],
        "local_id": "84",
        "full_desc": "<input bound_box=220,71,807,202>google.com.hk/search?gs_ssp=eJzj4tTP1TcwMU02T1JgNG</input>",
        "desc": "<input bound_box=220,71,807,202>google.com.hk/search?gs_ssp=eJzj4tTP1TcwMU02T1JgNG</input>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            683,
            684
        ],
        "focused": false,
        "bounds": [
            [
                828,
                63
            ],
            [
                1080,
                210
            ]
        ],
        "resource_id": "com.android.chrome:id/toolbar_buttons",
        "checked": false,
        "text": null,
        "class": "android.widget.LinearLayout",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 676,
        "temp_id": 682,
        "size": "252*147",
        "signature": "[class]android.widget.LinearLayout[resource_id]com.android.chrome:id/toolbar_buttons[visible]True[text]None[enabled,,]",
        "view_str": "e58903a2438d4a5dab10eda3de6ac2d7",
        "bound_box": "828,63,1080,210",
        "content_free_signature": "[class]android.widget.LinearLayout[resource_id]com.android.chrome:id/toolbar_buttons[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "3 open tabs, tap to switch tabs",
        "children": [],
        "focused": false,
        "bounds": [
            [
                828,
                63
            ],
            [
                954,
                210
            ]
        ],
        "resource_id": "com.android.chrome:id/tab_switcher_button",
        "checked": false,
        "text": null,
        "class": "android.widget.ImageButton",
        "scrollable": false,
        "selected": false,
        "long_clickable": true,
        "parent": 682,
        "temp_id": 683,
        "size": "126*147",
        "signature": "[class]android.widget.ImageButton[resource_id]com.android.chrome:id/tab_switcher_button[visible]True[text]None[enabled,,]",
        "view_str": "154aa901cf2539a34313cac7044838e7",
        "bound_box": "828,63,954,210",
        "content_free_signature": "[class]android.widget.ImageButton[resource_id]com.android.chrome:id/tab_switcher_button[visible]True",
        "allowed_actions": [
            "touch",
            "long_touch"
        ],
        "status": [],
        "local_id": "85",
        "full_desc": "<button alt='3 open tabs, tap to switch tabs' bound_box=828,63,954,210></button>",
        "desc": "<button alt='3 open tabs, tap to switch tabs' bound_box=828,63,954,210></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 2,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            685,
            686
        ],
        "focused": false,
        "bounds": [
            [
                954,
                63
            ],
            [
                1080,
                210
            ]
        ],
        "resource_id": "com.android.chrome:id/menu_button_wrapper",
        "checked": false,
        "text": null,
        "class": "android.widget.FrameLayout",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 682,
        "temp_id": 684,
        "size": "126*147",
        "signature": "[class]android.widget.FrameLayout[resource_id]com.android.chrome:id/menu_button_wrapper[visible]True[text]None[enabled,,]",
        "view_str": "1e1ead4d212396af21505c5794826e6a",
        "bound_box": "954,63,1080,210",
        "content_free_signature": "[class]android.widget.FrameLayout[resource_id]com.android.chrome:id/menu_button_wrapper[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": true,
        "is_password": false,
        "focusable": true,
        "enabled": true,
        "content_description": "Update available. More options",
        "children": [],
        "focused": false,
        "bounds": [
            [
                954,
                63
            ],
            [
                1080,
                210
            ]
        ],
        "resource_id": "com.android.chrome:id/menu_button",
        "checked": false,
        "text": null,
        "class": "android.widget.ImageButton",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 684,
        "temp_id": 685,
        "size": "126*147",
        "signature": "[class]android.widget.ImageButton[resource_id]com.android.chrome:id/menu_button[visible]True[text]None[enabled,,]",
        "view_str": "48d13517bb485302c3b98bb39ffc89d8",
        "bound_box": "954,63,1080,210",
        "content_free_signature": "[class]android.widget.ImageButton[resource_id]com.android.chrome:id/menu_button[visible]True",
        "allowed_actions": [
            "touch"
        ],
        "status": [],
        "local_id": "86",
        "full_desc": "<button alt='Update available. More options' bound_box=954,63,1080,210></button>",
        "desc": "<button alt='Update available. More options' bound_box=954,63,1080,210></button>"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                954,
                63
            ],
            [
                1080,
                210
            ]
        ],
        "resource_id": "com.android.chrome:id/menu_badge",
        "checked": false,
        "text": null,
        "class": "android.widget.ImageView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 684,
        "temp_id": 686,
        "size": "126*147",
        "signature": "[class]android.widget.ImageView[resource_id]com.android.chrome:id/menu_badge[visible]True[text]None[enabled,,]",
        "view_str": "26549dd4b1f649a3d7fe770605c574d7",
        "bound_box": "954,63,1080,210",
        "content_free_signature": "[class]android.widget.ImageView[resource_id]com.android.chrome:id/menu_badge[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": true,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                210
            ],
            [
                1080,
                231
            ]
        ],
        "resource_id": "com.android.chrome:id/toolbar_shadow",
        "checked": false,
        "text": null,
        "class": "android.widget.ImageView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 675,
        "temp_id": 687,
        "size": "1080*21",
        "signature": "[class]android.widget.ImageView[resource_id]com.android.chrome:id/toolbar_shadow[visible]True[text]None[enabled,,]",
        "view_str": "4231d165ebbf1f8ff621fd38bc114f6f",
        "bound_box": "0,210,1080,231",
        "content_free_signature": "[class]android.widget.ImageView[resource_id]com.android.chrome:id/toolbar_shadow[visible]True"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                1,
                205
            ],
            [
                1,
                210
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.widget.ImageView",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 674,
        "temp_id": 688,
        "size": "0*5",
        "signature": "[class]android.widget.ImageView[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "0a712eaeb10310c39b221526856e512e",
        "bound_box": "1,205,1,210",
        "content_free_signature": "[class]android.widget.ImageView[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            690
        ],
        "focused": false,
        "bounds": [
            [
                0,
                2274
            ],
            [
                1080,
                2274
            ]
        ],
        "resource_id": "com.android.chrome:id/bottom_container",
        "checked": false,
        "text": null,
        "class": "android.widget.FrameLayout",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 5,
        "temp_id": 689,
        "size": "1080*0",
        "signature": "[class]android.widget.FrameLayout[resource_id]com.android.chrome:id/bottom_container[visible]False[text]None[enabled,,]",
        "view_str": "85eac73d1925c7ff6cae83a28573f164",
        "bound_box": "0,2274,1080,2274",
        "content_free_signature": "[class]android.widget.FrameLayout[resource_id]com.android.chrome:id/bottom_container[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 1,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [
            691
        ],
        "focused": false,
        "bounds": [
            [
                0,
                2274
            ],
            [
                1080,
                2274
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.widget.FrameLayout",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 689,
        "temp_id": 690,
        "size": "1080*0",
        "signature": "[class]android.widget.FrameLayout[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "e52539f6dce797acd524467109d49286",
        "bound_box": "0,2274,1080,2274",
        "content_free_signature": "[class]android.widget.FrameLayout[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                2274
            ],
            [
                1080,
                2274
            ]
        ],
        "resource_id": null,
        "checked": false,
        "text": null,
        "class": "android.widget.FrameLayout",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 690,
        "temp_id": 691,
        "size": "1080*0",
        "signature": "[class]android.widget.FrameLayout[resource_id]None[visible]False[text]None[enabled,,]",
        "view_str": "e9f953084c0e6f3b3f412cd2cd2ce4c3",
        "bound_box": "0,2274,1080,2274",
        "content_free_signature": "[class]android.widget.FrameLayout[resource_id]None[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                2274
            ],
            [
                1080,
                2274
            ]
        ],
        "resource_id": "com.android.chrome:id/navigation_popup_anchor_stub",
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 4,
        "temp_id": 692,
        "size": "1080*0",
        "signature": "[class]android.view.View[resource_id]com.android.chrome:id/navigation_popup_anchor_stub[visible]False[text]None[enabled,,]",
        "view_str": "77afc2be9104e5b04d71a00d961bb848",
        "bound_box": "0,2274,1080,2274",
        "content_free_signature": "[class]android.view.View[resource_id]com.android.chrome:id/navigation_popup_anchor_stub[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                2274
            ],
            [
                0,
                2274
            ]
        ],
        "resource_id": "com.android.chrome:id/menu_anchor_stub",
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 4,
        "temp_id": 693,
        "size": "0*0",
        "signature": "[class]android.view.View[resource_id]com.android.chrome:id/menu_anchor_stub[visible]False[text]None[enabled,,]",
        "view_str": "85dac7e76bd588b46f4fb99022c9bac9",
        "bound_box": "0,2274,0,2274",
        "content_free_signature": "[class]android.view.View[resource_id]com.android.chrome:id/menu_anchor_stub[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                0
            ],
            [
                1080,
                63
            ]
        ],
        "resource_id": "android:id/statusBarBackground",
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 0,
        "temp_id": 694,
        "size": "1080*63",
        "signature": "[class]android.view.View[resource_id]android:id/statusBarBackground[visible]False[text]None[enabled,,]",
        "view_str": "e521e91baefa4fd89e4dc021110f2ae7",
        "bound_box": "0,0,1080,63",
        "content_free_signature": "[class]android.view.View[resource_id]android:id/statusBarBackground[visible]False"
    },
    {
        "package": "com.android.chrome",
        "visible": false,
        "checkable": false,
        "child_count": 0,
        "editable": false,
        "clickable": false,
        "is_password": false,
        "focusable": false,
        "enabled": true,
        "content_description": null,
        "children": [],
        "focused": false,
        "bounds": [
            [
                0,
                2274
            ],
            [
                1080,
                2400
            ]
        ],
        "resource_id": "android:id/navigationBarBackground",
        "checked": false,
        "text": null,
        "class": "android.view.View",
        "scrollable": false,
        "selected": false,
        "long_clickable": false,
        "parent": 0,
        "temp_id": 695,
        "size": "1080*126",
        "signature": "[class]android.view.View[resource_id]android:id/navigationBarBackground[visible]False[text]None[enabled,,]",
        "view_str": "ad4baa7317b83af5de62c848ffcc94cf",
        "bound_box": "0,2274,1080,2400",
        "content_free_signature": "[class]android.view.View[resource_id]android:id/navigationBarBackground[visible]False"
    }
]